`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,
	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:12] == 4'b1011);	// B000-B001 : KIA (B002-BFFF = repeats)
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)};
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h0000000000000F001E160A01647257051001210A10016F6C4805102A03000000,
progmem.ram00.INIT_01 = 256'h666006667E787C3C2004003C1C0C3C180000000C381866000000000000000000,
progmem.ram00.INIT_02 = 256'h000000FF020820803618000000080000001800601C06603018007E66C67E7C7C,
progmem.ram00.INIT_03 = 256'h102010202E281020C03038007C08381038003828100010000000FF8080E0FFFF,
progmem.ram00.INIT_04 = 256'h0000000000000F00402808022810204810201020002810102028083C28102070,
progmem.ram00.INIT_05 = 256'h76600666606C6666300C1866301C6624000024186C3E66000000000000000000,
progmem.ram00.INIT_06 = 256'h00000000020820806C18000000180000001818603006601818600666C6186666,
progmem.ram00.INIT_07 = 256'h281028105800281020104400F410042874001C001044380000007FC040E0FFFF,
progmem.ram00.INIT_08 = 256'h0000000000000F004000103C0028103028102810000028082000104C00281048,
progmem.ram00.INIT_09 = 256'h766006666066666E18181866603C066600001830685824000000000000000000,
progmem.ram00.INIT_0A = 256'h0000FF000208208000187E66663C5E7C5C18007C303E7C0C3C300C3C6C186666,
progmem.ram00.INIT_0B = 256'h38387C7C58000000C4104400F40018106C7C64001038540007E03FE020E0FF00,
progmem.ram00.INIT_0C = 256'h0000000000000F005844444C38383808000038386C3838383800005438383844,
progmem.ram00.INIT_0D = 256'h7E60067E78667C6A0C30003C7C6C0C6600007E30323C00000000000000000000,
progmem.ram00.INIT_0E = 256'h000000000208208000180C3C66186066661818667C6666003C1818186C187C7C,
progmem.ram00.INIT_0F = 256'h101040408C101010287C38007400200074043C000028500018181FF010E0FF00,
progmem.ram00.INIT_10 = 256'h00000000000F00006444445444444438303044441204040424444454444444E4,
progmem.ram00.INIT_11 = 256'h6E6066666066666618180066667E3066001018306C1A00000000000000000000,
progmem.ram00.INIT_12 = 256'h00FF000002082080001818183C1860666618186630666600660C303C38187860,
progmem.ram00.INIT_13 = 256'h10106070F8282828D408000014003C006C007C001038540010080FF808E00000,
progmem.ram00.INIT_14 = 256'h00000000000F0000644444644444444410107C7C7E3C3C3C3844445444444444,
progmem.ram00.INIT_15 = 256'h6E606666606C6660300C1866660C6024181824186C7C00000000000000000000,
progmem.ram00.INIT_16 = 256'h00000000020820800018303C3C18607C66181866306666000006606638186C60,
progmem.ram00.INIT_17 = 256'h10104040884444442C287C00140000006C00000010443800200407FC04E00000,
progmem.ram00.INIT_18 = 256'h00000000000F0000584444784444444410104040904444442044446444444448,
progmem.ram00.INIT_19 = 256'h667E3C6660787C3C2004183C3C0C7E181810000C3A1800000000000000000000,
progmem.ram00.INIT_1A = 256'hFF0000000208208000187E66180C6060660C1866303E7C0000007E6610186660,
progmem.ram00.INIT_1B = 256'h38387C7C8E7C7C7C5C380008140000003800000010001000200403FE02E00000,
progmem.ram00.INIT_1C = 256'h00000000000F00004038388038383838383838386E3C3C3C2038387838383870,
progmem.ram00.INIT_1D = 256'h0000000000000000000000000000000000200000000000000000000000000000,
progmem.ram00.INIT_1E = 256'h0000000002082080000000000000006000007000000000000000000000000000,
progmem.ram00.INIT_1F = 256'h000000000044444404080010000000000000000000000000200401FF01E00000,
progmem.ram00.INIT_20 = 256'h10A030C050E07000400000000000000000000000000000000000000000000000,
progmem.ram00.INIT_21 = 256'h6400237400006AE06A0000000000000000000000000070009020B040D060F080,
progmem.ram00.INIT_22 = 256'h0000A8E030425E5E12A800008EE0940076A0E0A464178E000000746412026414,
progmem.ram00.INIT_23 = 256'h001366126466A1EC000000D86612306814D80000BC2E640041015C16AAC8E0BC,
progmem.ram00.INIT_24 = 256'h42E0EE3CE0EE36E0EE30E0DA2AE0006860A1BE1CE010000000EC641250641466,
progmem.ram00.INIT_25 = 256'h5EE05C01135C6012016014126AE05E000010E0EE5AE0EE54E0EE4EE0EE48E0EE,
progmem.ram00.INIT_26 = 256'hAAE090BCE0640030AA000000805C503100806212FF62146092E0A06217800000,
progmem.ram00.INIT_27 = 256'hE200E00200F00000E02E5A5A41E00000C0E0C60082D8E0DC0017B05C14C00000,
progmem.ram00.INIT_28 = 256'h285A31045A141A34E0280000182E035A1418000004E0E214E00600040000F0E0,
progmem.ram00.INIT_29 = 256'h702E025A14700000602E025A14600000502E015A1450000000425AA142000000,
progmem.ram00.INIT_2A = 256'h5C0062BCE0B00000A02E065A14A0000090E0529CE0900000802E045A14800000,
progmem.ram00.INIT_2B = 256'h5E0052FCE05C0062F2E0E60000B0E0C2E2E06004135A62121AD0E05E0052C6E0,
progmem.ram00.INIT_2C = 256'hE04210174438E0480000B0156228E01C0000E6E06C18E06004135A62121A06E0,
progmem.ram00.INIT_2D = 256'h00004CE0E878E04CE07211174468E0780000D8156258E04C00001CE0B248E01C,
progmem.ram00.INIT_2E = 256'hBA0000B0E0B0000086E006ACE086E0F2A2E0A60040F0164492E08600007CE07C,
progmem.ram00.INIT_2F = 256'hE0F80000EEE0EE0000BAE0E2EAE00800B2E0E0BAE088D6E0DA0030F01644C6E0,
progmem.ram00.INIT_30 = 256'h15523EE054001A34E0280000F8E00624E0F01EE0F8E0BC14E0180020F0164404,
progmem.ram00.INIT_31 = 256'hE02A7EE058E0FA74E0780010F0164464E058000028E04E54E01E4EE0540000EE,
progmem.ram00.INIT_32 = 256'h01C610015A15AE000088E0F2AAE088E05AA0E0A400174494E088000058E02A84,
progmem.ram00.INIT_33 = 256'h0642F60000CAE0F2F2E0D0008AE8E0EC011744DCE0B0D6E0CA0000AEE0E2C6E0,
progmem.ram00.INIT_34 = 256'h41FF54160156142C000010E0CC28E0F822E0AC1CE0100000F62E5A2156561202,
progmem.ram00.INIT_35 = 256'h007056003170000056E0560056FF246C56175600002CE0005656410152710001,
progmem.ram00.INIT_36 = 256'h16B8000094E012B4E082AEE00094A81201581694000000805612FF5414800000,
progmem.ram00.INIT_37 = 256'hDCE012FCE02EF6E000DCF0127A5816DC0000B8E012D8E072D2E000B8CC126C58,
progmem.ram00.INIT_38 = 256'h58021334000024E054061324000000E01220E0581AE0000014127D5816000000,
progmem.ram00.INIT_39 = 256'h7A000064E06A761E01001564000048E002521B58581200021648000000340212,
progmem.ram00.INIT_3A = 256'hE0C800E0021666B4E0A800007AE04AA4E0669EE002007AE03690E09400F00216,
progmem.ram00.INIT_3B = 256'h00D2E0D80096F6E0BAF0E0DEEAE002E4E0AADEE0D20000A8E0AE021EA8E07CC4,
progmem.ram00.INIT_3C = 256'h00000000000000000000000000000000FEE0D41CE01216E07210E0260AE0FE00,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'h00000000000F00F000000000216C6F06060021020500006C6505050000000F1E,
progmem.ram01.INIT_01 = 256'h3C42663C3C7E1E103C00003C7E7E3C080000003018706C180000000000000000,
progmem.ram01.INIT_02 = 256'h0000000001041040AA300C00000000000000600000000000003C3C6666663C3C,
progmem.ram01.INIT_03 = 256'h280828083810340810300010000038107C000038384418102004FF0101F0C0FF,
progmem.ram01.INIT_04 = 256'h00000000000F00F0280810200034083428082808001034083008102000340834,
progmem.ram01.INIT_05 = 256'h66666C186060303866001866064066180600181818546C180000000000000000,
progmem.ram01.INIT_06 = 256'h000000FF0104104055181800000000000000601800000000000C306666666666,
progmem.ram01.INIT_07 = 256'h0010001044285810001050300000041000001454404420002004FE0302F0C0FF,
progmem.ram01.INIT_08 = 256'h00000000000F00F0001028101058105800100010002858104810281044581058,
progmem.ram01.INIT_09 = 256'h667E781860606038067E18660C7C06380C00180C1868FE180000000000000000,
progmem.ram01.INIT_0A = 256'h0000000001041040AA181866C6663E3E3CFC66003E3C3E3C000C303C66666066,
progmem.ram01.INIT_0B = 256'h38387C7C401000001010281000441C7C0000286C382820102004FC0704F0C0FF,
progmem.ram01.INIT_0C = 256'h00000000000F00F0444400440038385800003838381038385044000028383844,
progmem.ram01.INIT_0D = 256'h667E70186E78606C0C00003E0C061C18187E7E0C00106C180000000000000000,
progmem.ram01.INIT_0E = 256'h0000FF000104104055066066C666606666D66C3866666006000C303C7E663C66,
progmem.ram01.INIT_0F = 256'h1010404040101010207C14101044041000385064447C70101008F80F08F0C000,
progmem.ram01.INIT_10 = 256'h0000000000F0F000444444447C44446430304444443804047828444410444464,
progmem.ram01.INIT_11 = 256'h666678186660607C187E1806180606183000180C002CFE180000000000000000,
progmem.ram01.INIT_12 = 256'h0000000001041040AA181866D6663C6666D67818667E603E000C30187E660666,
progmem.ram01.INIT_13 = 256'h101070704028282840302810004438100000286C381020101818F01F10F0C000,
progmem.ram01.INIT_14 = 256'h0000000000F0F000444444440044444410107C7C401C3C3C4410444428444454,
progmem.ram01.INIT_15 = 256'h66666C18666030C60000180C186666186000181800546C000000000000000000,
progmem.ram01.INIT_16 = 256'h00FF0000010410405518183ED666063E66C66C183E606066000C30186666666E,
progmem.ram01.INIT_17 = 256'h1010404044444444440850000064000000001454047C201007E0E03F20F0C000,
progmem.ram01.INIT_18 = 256'h0000000000F0F0003C3C4444104444441010404044644444641044444444444C,
progmem.ram01.INIT_19 = 256'h3C66663C3C7E1EC618001038183C3C3C00000030001C6C180000000000000000,
progmem.ram01.INIT_1A = 256'h0000000001041040AA300C067C3A7C063CC6663C063C3E3A7E3C3C18423C3C3C,
progmem.ram01.INIT_1B = 256'h38387C7C387C7C7C38100000005C007C0000003838105C100000C07F40F0C000,
progmem.ram01.INIT_1C = 256'h0000000000F0F000040438380038384438383838383C3C3C5810383800383844,
progmem.ram01.INIT_1D = 256'h0000000000000000000020000000000000000000000000000000000000000000,
progmem.ram01.INIT_1E = 256'hFF000000010410405500003C00000006000000003C0000000000000000000006,
progmem.ram01.INIT_1F = 256'h000000006044444400380000004000000000000000000000000080FF80F0C000,
progmem.ram01.INIT_20 = 256'h1814110D0A060300383800000000000000000000600000008000000000000000,
progmem.ram01.INIT_21 = 256'h080011081300081208130000000000000000000000003A3733302C2925221E1B,
progmem.ram01.INIT_22 = 256'h1300081208410808120813000812081E080811080812081300E0080813000812,
progmem.ram01.INIT_23 = 256'h0114082B080812081300E008081300081A081300083108C04100081208081108,
progmem.ram01.INIT_24 = 256'h091108091108091108091108091130080812080911091300E008081300081208,
progmem.ram01.INIT_25 = 256'h0912080014080813000812090911091300091208091108091108091108091108,
progmem.ram01.INIT_26 = 256'h091208091108C0110913002E09080011E0090813FF0812090911090812091300,
progmem.ram01.INIT_27 = 256'h090A11001009130009310808120913000912091E090911098015FF0812091300,
progmem.ram01.INIT_28 = 256'h0A08410008120A0A110A13000AA10008120A13000A12090A1100100A13000912,
progmem.ram01.INIT_29 = 256'h0A210008120A13000AA10008120A13000AA10008120A13002E0A08120A13002E,
progmem.ram01.INIT_2A = 256'h08130A0A110A13000AA10008120A13000A120A0A110A13000A210008120A1300,
progmem.ram01.INIT_2B = 256'h08130A0A1108130A0A110A13000A12090A110800140808130A0A1108130A0A11,
progmem.ram01.INIT_2C = 256'h120B00160A0B110B1780FF140A0B110B13000A12080B110800140808130A0B11,
progmem.ram01.INIT_2D = 256'h13000B120A0B110B120B00160A0B110B1780FF140A0B110B13000B120A0B110B,
progmem.ram01.INIT_2E = 256'h0B13000B120B13000B120A0B110B12090B110B170000150A0B110B13000B120B,
progmem.ram01.INIT_2F = 256'h110B13000B120B13000B12090B1100100B0B110B120B0B110B170000150A0B11,
progmem.ram01.INIT_30 = 256'h140A0C110C170A0C110C13000B120A0C110B0C110B120B0C110C170000150A0C,
progmem.ram01.INIT_31 = 256'h110C0C110C120B0C110C170000150A0C110C13000C120B0C110B0C110C1780FF,
progmem.ram01.INIT_32 = 256'h000C170008120C13000C12090C110C120C0C110C00160A0C110C13000C120A0C,
progmem.ram01.INIT_33 = 256'h00110C13000C12090C110C1E0C0C110C00160A0C110C0C110C13000C12090C11,
progmem.ram01.INIT_34 = 256'h14FF08120008120D13000D120C0D110C0D11090D110D13000C31084408081200,
progmem.ram01.INIT_35 = 256'h2E0D0800110D13000D12081308FF110D08120D13000D1230080812000D518000,
progmem.ram01.INIT_36 = 256'h120D13000D120D0D110D0D11E00D0D170008120D1300E00D0813FF08120D1300,
progmem.ram01.INIT_37 = 256'h0D120D0D110D0D11E00D0D170008120D13000D120D0D110D0D11E00D0D170008,
progmem.ram01.INIT_38 = 256'h08B01A0E13000E120800120E13000E120D0E110D0E11E00E0E170008120E1300,
progmem.ram01.INIT_39 = 256'h0E13000E120E0E1700B01A0E13000E12B0C01308081380B01A0E1300E00EB01B,
progmem.ram01.INIT_3A = 256'h110E1700B01A0E0E110E13000E120E0E110E0E11B01B0E120E0E110E1700B01A,
progmem.ram01.INIT_3B = 256'h000E120E1E0D0E110D0E110D0E110E0E110E0E110E13000E120EB01B0E120E0E,
progmem.ram01.INIT_3C = 256'h000000000000000000000000000000000E120E0F110D0F110D0F110E0F110E13,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
