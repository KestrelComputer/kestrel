`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:		12:51:57 11/06/2011 
// Design Name:		Kestrel-2 rev 1A
// Module Name:		M_kestrel2 
// Project Name:		Kestrel-2
// Target Devices:	NEXYS2
// Tool versions: 
// Description: 
//		The Kestrel 2 computer, top-level integration module.
//
// Dependencies: 
//		M_uxa, M_mem, M_j1a
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module M_kestrel2(
	output N2_CA_O,
	output N2_CB_O,
	output N2_CC_O,
	output N2_CD_O,
	output N2_CE_O,
	output N2_CF_O,
	output N2_CG_O,
	output N2_DP_O,
	output N2_A0_O,
	output N2_A1_O,
	output N2_A2_O,
	output N2_A3_O,
	output N2_HSYNC_O,
	output N2_VSYNC_O,
	output [2:0] N2_RED_O,
	output [2:0] N2_GRN_O,
	output [2:1] N2_BLU_O,
	input N2_PS2D_I,
	input N2_PS2C_I,
	input N2_50MHZ_I,
	input N2_RST_I
);

	// Permanently hold the LED outputs in an inactive state,
	// to prevent unnecessary current draw on the part of the
	// FPGA.
	reg a_, b_, c_, d_, e_, f_, g_, dp_, a0_, a1_, a2_, a3_;
	assign N2_CA_O = a_;
	assign N2_CB_O = b_;
	assign N2_CC_O = c_;
	assign N2_CD_O = d_;
	assign N2_CE_O = e_;
	assign N2_CF_O = f_;
	assign N2_CG_O = g_;
	assign N2_DP_O = dp_;
	assign N2_A0_O = a0_;
	assign N2_A1_O = a1_;
	assign N2_A2_O = a2_;
	assign N2_A3_O = a3_;

	initial begin
		a_ <= 1;		e_ <= 1;
		b_ <= 1;		f_ <= 1;
		c_ <= 1;		g_ <= 1;
		d_ <= 1;		dp_ <= 1;
		a0_ <= 1; 	a1_ <= 1;
		a2_ <= 1; 	a3_ <= 1;
	end

	// Each major module has its own set of inputs and
	// outputs.  We declare them here so that the synthesizer
	// has complete knowledge of what to expect before we start
	// routing signals around.
	wire [13:1] j1a_ins_adr_o;
	wire [15:0] j1a_ins_dat_i;
	wire        j1a_ins_cyc_o;
	wire [15:1] j1a_dat_adr_o;
	reg  [15:0] j1a_dat_dat_i;
	wire [15:0] j1a_dat_dat_o;
	wire        j1a_dat_cyc_o;
	wire        j1a_dat_we_o;
	wire        j1a_stb_o;
	reg         j1a_ack_i;

	wire			pm_dat_ack_o;
	wire			pm_ins_ack_o;
	wire [15:0]	pm_dat_o;
	reg 			pm_dat_stb;

	wire [15:0]	vm_dat_o;
	reg			vm_dat_stb;
	wire			vm_dat_ack_o;

	wire [13:1]	mgia_adr_o;
	wire [15:0]	mgia_dat_i;
	wire			mgia_cyc_o;
	wire			mgia_stb_o;
	wire			mgia_ack_i;
	wire			sys_clk;

	// Instantiate the J1A microprocessor.
	M_j1a j1a(
		.sys_res_i(N2_RST_I),
		.sys_clk_i(sys_clk),
		.ins_adr_o(j1a_ins_adr_o),
		.ins_dat_i(j1a_ins_dat_i),
		.dat_adr_o(j1a_dat_adr_o),
		.dat_dat_o(j1a_dat_dat_o),
		.dat_dat_i(j1a_dat_dat_i),
		.dat_we_o(j1a_dat_we_o),
		.dat_cyc_o(j1a_dat_cyc_o),
		.ins_cyc_o(j1a_ins_cyc_o),
		.shr_stb_o(j1a_stb_o),
		.shr_ack_i(j1a_ack_i)
	);

	wire data_access = ~N2_RST_I & j1a_stb_o & j1a_dat_cyc_o;
	wire addressing_prg_mem = j1a_dat_adr_o[15:14] == 2'b00;
	wire addressing_vid_mem = j1a_dat_adr_o[15:14] == 2'b10;

	always @* begin
		// When fetching data from various resources, the CPU will
		// need to select which output data bus to read from.
		if (addressing_prg_mem)
			j1a_dat_dat_i <= pm_dat_o;
		else if (addressing_vid_mem)
			j1a_dat_dat_i <= vm_dat_o;
//		else if (addressing_kbd_ps2)
//			j1a_dat_dat_i <= kbd_dat_o;
		else
			j1a_dat_dat_i <= 16'hxxxx;
			
		// Peripherals won't know to drive their buses, however,
		// unless told to do so by asserting the appropriate
		// data strobes.
		pm_dat_stb <= data_access & addressing_prg_mem;
		vm_dat_stb <= data_access & addressing_vid_mem;

		// Since the Kestrel-2 lacks multi-master support,
		// we can get by with simply ORing all the acknowledgements
		// together.
		j1a_ack_i <= pm_ins_ack_o | pm_dat_ack_o | vm_dat_ack_o;
	end

	// Program Memory ($0000-$3FFF)
	M_mem pm(
		.ins_adr_i(j1a_ins_adr_o),
		.ins_dat_o(j1a_ins_dat_i),
		.ins_cyc_i(j1a_ins_cyc_o),
		.ins_stb_i(j1a_stb_o),
		.ins_ack_o(pm_ins_ack_o),

		.dat_adr_i(j1a_dat_adr_o[13:1]),
		.dat_dat_o(pm_dat_o),
		.dat_dat_i(j1a_dat_dat_o),
		.dat_we_i(j1a_dat_we_o),
		.dat_cyc_i(j1a_dat_cyc_o),
		.dat_stb_i(pm_dat_stb),
		.dat_ack_o(pm_dat_ack_o),

		.sys_clk_i(sys_clk),
		.sys_rst_i(N2_RST_I)
	);
	
	// Video Memory ($8000-$BFFF)
	M_mem vm(
		.ins_adr_i(mgia_adr_o),
		.ins_dat_o(mgia_dat_i),
		.ins_cyc_i(mgia_cyc_o),
		.ins_stb_i(mgia_stb_o),
		.ins_ack_o(mgia_ack_i),
		
		.dat_adr_i(j1a_dat_adr_o[13:1]),
		.dat_dat_o(vm_dat_o),
		.dat_dat_i(j1a_dat_dat_o),
		.dat_we_i(j1a_dat_we_o),
		.dat_cyc_i(j1a_dat_cyc_o),
		.dat_stb_i(vm_dat_stb),
		.dat_ack_o(vm_dat_ack_o),
		
		.sys_clk_i(sys_clk),
		.sys_rst_i(N2_RST_I)
	);

	// Monochrome Graphics Interface Adapter
	M_uxa_mgia mgia(
		.CLK_I_50MHZ(N2_50MHZ_I),
		.RST_I(N2_RST_I),
		.CLK_O_25MHZ(sys_clk),

		.HSYNC_O(N2_HSYNC_O),
		.VSYNC_O(N2_VSYNC_O),
		.RED_O(N2_RED_O),
		.GRN_O(N2_GRN_O),
		.BLU_O(N2_BLU_O),
	
		.MGIA_ADR_O(mgia_adr_o),
		.MGIA_DAT_I(mgia_dat_i),
		.MGIA_CYC_O(mgia_cyc_o),
		.MGIA_STB_O(mgia_stb_o),
		.MGIA_ACK_I(mgia_ack_i)
	);

	// Keyboard PS2IO ($FFFE)
	
	// Video RAM static image (at boot-time)
	defparam
vm.ram00_07.INIT_3F = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_3E = 256'h55555555555555555555555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_3D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_3C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_3B = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_3A = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_39 = 256'h55555555555555555555000000000000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_38 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_37 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA000C228AF1C2,
vm.ram00_07.INIT_36 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_35 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_34 = 256'h55555555555555555555010C228A8882AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_33 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_32 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA019822FA8882,
vm.ram00_07.INIT_31 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_30 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_2F = 256'h55555555555555555555C1D82A53F082AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_2E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_2D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA21F02A528882,
vm.ram00_07.INIT_2C = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_2B = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_2A = 256'h5555555555555555555521FC36228882AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_29 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_28 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAC1F8A223F1CF,
vm.ram00_07.INIT_27 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_26 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_25 = 256'h5555555555555555555501F000000000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_24 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_23 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAE1E0A0FB7228,
vm.ram00_07.INIT_22 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_21 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_20 = 256'h5555555555555555555501C0A0828A28AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_1F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_1E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA0180A0820A28,
vm.ram00_07.INIT_1D = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_1C = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_1B = 256'h555555555555555555558100BC8373EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_1A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_19 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA0000A282822A,
vm.ram00_07.INIT_18 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_17 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_16 = 256'h555555555555555555550000A282894DAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_15 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_14 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAE000BC837088,
vm.ram00_07.INIT_13 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_12 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_11 = 256'h55555555555555555555000000000000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_10 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_0F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAEF88088B8BE7,
vm.ram00_07.INIT_0E = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_0D = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_0C = 256'h55555555555555555555080088929208AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_0B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_0A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA080888A2A200,
vm.ram00_07.INIT_09 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_08 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_07 = 256'h55555555555555555555880808F3C387AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_06 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_05 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA081C088AA208,
vm.ram00_07.INIT_04 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_03 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
vm.ram00_07.INIT_02 = 256'h55555555555555555555081C888A9208AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_01 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
vm.ram00_07.INIT_00 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAE8083EF38BE7;

	// System Firmware


defparam
    pm.ram00_07.INIT_00 = 256'h6181710F710F6180200E4001620380016203660061816181730F6600FFFF125E,
    pm.ram00_07.INIT_01 = 256'h401A20226303800160817C0C710F6180710F2018400162038001620366006181,
    pm.ram00_07.INIT_02 = 256'h61806403630380FF401A61816D0380086180730F80FF69038008401A730F80FF,
    pm.ram00_07.INIT_03 = 256'h80016081710F6123618064036303660080FF401A6181630380FF6180710F6123,
    pm.ram00_07.INIT_04 = 256'h7D0F80047D0F8003710F6103612361806203401A618161810027003220436303,
    pm.ram00_07.INIT_05 = 256'h0000700C80BE0000700C80B8004C40507D0F8008720F6D03800260816D038004,
    pm.ram00_07.INIT_06 = 256'h00000000000000000000000F0F0000F0700C80D00000700C80CA0000700C80C4,
    pm.ram00_07.INIT_07 = 256'h0000000000000C3038181870666C001800000000000000000000000000000000,
    pm.ram00_07.INIT_08 = 256'h663C60420666663C7E3C787E7C1E3C10203C040000003C3C1C7E0C7E3C3C1808,
    pm.ram00_07.INIT_09 = 256'h00001800006060001C000600600030001800003C7E3C6666C6667E667C3C7C3C,
    pm.ram00_07.INIT_0A = 256'h000000000000FF00020108042010804036AA1830000C00000000080000000000,
    pm.ram00_07.INIT_0B = 256'h387C000038002838103800441018001000200004FFFF80018001E0F0FFC0FFFF,
    pm.ram00_07.INIT_0C = 256'h10282008102820082E38281010342008C0103030380000107C00080038381010,
    pm.ram00_07.INIT_0D = 256'h102820081028200800002810103410082030280808103C202800103420087034,
    pm.ram00_07.INIT_0E = 256'h00000000000000000000000F0F0000F040282808081002202800103420084834,
    pm.ram00_07.INIT_0F = 256'h00060000241818186C183E54666C001800000000000000000000000000000000,
    pm.ram00_07.INIT_10 = 256'h76666066066C661860606C606630663830660C001818666630061C4066662418,
    pm.ram00_07.INIT_11 = 256'h000018001860601830000600600018001800600C06306666C666186666666666,
    pm.ram00_07.INIT_12 = 256'h00000000000000FF02010804201080406C551818001800000000180000000000,
    pm.ram00_07.INIT_13 = 256'h740000001C1400541040444438200000002000047FFEC0034002E0F0FFC0FFFF,
    pm.ram00_07.INIT_14 = 256'h280010102800101058440028285810102000101044500030F400100004042810,
    pm.ram00_07.INIT_15 = 256'h280010102800101000000028285808102048001010284C100044285810104858,
    pm.ram00_07.INIT_16 = 256'h00000000000000000000000F0F0000F04000001010283C100010285810103058,
    pm.ram00_07.INIT_17 = 256'h000C00001818300C6818586824FE001800000000000000000000000000000000,
    pm.ram00_07.INIT_18 = 256'h7666607E067866186060666066606E381806187E18186666600C3C7C06066638,
    pm.ram00_07.INIT_19 = 256'h5C3C18FC00667C00303E3E3C7C3E0C3C3C00300C0C303C3C6C66186666606666,
    pm.ram00_07.INIT_1A = 256'h00000000FF000000020108042010804000AA18187E18666666C63C665E3E7C3E,
    pm.ram00_07.INIT_1B = 256'h6C007C006428006C10383828542000100720E0043FFCE0072004E0F0FFC000FF,
    pm.ram00_07.INIT_1C = 256'h383838387C7C7C7C5840001000000000C410101044280010F4000044181C107C,
    pm.ram00_07.INIT_1D = 256'h00000000383838386C3838103838383838500044000054003828383838384444,
    pm.ram00_07.INIT_1E = 256'h00000000000000000000000F0F0000F05844444444004C443800383838380858,
    pm.ram00_07.INIT_1F = 256'h0018007E7E7E300C32003C10006C001800000000000000000000000000000000,
    pm.ram00_07.INIT_20 = 256'h7E66607E06707E18786E66787C606A6C0C0C300000003C3E7C0C6C060C1C6618,
    pm.ram00_07.INIT_21 = 256'h666618D6186C66387C666666666000063C00180C1830183C6C7E18667C3C7C66,
    pm.ram00_07.INIT_22 = 256'h0000000000FF00000201080420108040005518060C603C6666C6186660606666,
    pm.ram00_07.INIT_23 = 256'h740004383C5000640044287C50700010181018081FF8F00F1008E0F0FFC00000,
    pm.ram00_07.INIT_24 = 256'h10101010404040408C4010101010101028207C7C381400107410004420040010,
    pm.ram00_07.INIT_25 = 256'h303030304444444412440438040404042478442844445444441044444444E464,
    pm.ram00_07.INIT_26 = 256'h000000000000000000000FF000F000006444444444445444447C444444443864,
    pm.ram00_07.INIT_27 = 256'h003010001818300C6C001A2C00FE001800000000000000000000000000000000,
    pm.ram00_07.INIT_28 = 256'h6E66606666786618606666606660667C1818187E0018660666187E0630066618,
    pm.ram00_07.INIT_29 = 256'h666618D6187866183066667E6660003E66000C0C30303C18387E186678066066,
    pm.ram00_07.INIT_2A = 256'h0000FF0000000000020108042010804000AA1818181818663CD61866603C6666,
    pm.ram00_07.INIT_2B = 256'h6C0000007C28006C1038381054200010101808180FF0F81F0810E0F000C00000,
    pm.ram00_07.INIT_2C = 256'h1010101060707070F840282828282828D440083000280010140000443C380010,
    pm.ram00_07.INIT_2D = 256'h101010107C7C7C7C7E403C1C3C3C3C3C38444410444454444428444444444454,
    pm.ram00_07.INIT_2E = 256'h000000000000000000000FF000F0000064444444444464444400444444444444,
    pm.ram00_07.INIT_2F = 256'h18601800241818186C007C54006C000000000000000000000000000000000000,
    pm.ram00_07.INIT_30 = 256'h6E666066666C661860666C60663060C630000C001818660C66180C6660662418,
    pm.ram00_07.INIT_31 = 256'h666618C6186C6618303E6660666000660000060C60306618386618666C66606E,
    pm.ram00_07.INIT_32 = 256'h000000FF0000000002010804201080400055181830183C3E3CD6186660067C3E,
    pm.ram00_07.INIT_33 = 256'h6C000000001400541004447C38200010200704E007E0FC3F0420E0F000C00000,
    pm.ram00_07.INIT_34 = 256'h101010104040404088444444444444442C4428087C5000001400006400000000,
    pm.ram00_07.INIT_35 = 256'h101010104040404090444464444444442064441044446444444444444444484C,
    pm.ram00_07.INIT_36 = 256'h000000000000000000000FF000F00000583C443C444478444410444444444444,
    pm.ram00_07.INIT_37 = 256'h1800100000000C303A00181C006C001800000000000000000000000000000000,
    pm.ram00_07.INIT_38 = 256'h663C7E663C66663C603C787E7C1E3CC62018040018103C383C180C3C7E3C183C,
    pm.ram00_07.INIT_39 = 256'h663C0CC61866663C30063E3C7C3E003A007E003C7E3C66181042183C663C603C,
    pm.ram00_07.INIT_3A = 256'hFF00000000000000020108042010804000AA18307E0C6606187C0C3A607C6006,
    pm.ram00_07.INIT_3B = 256'h380000000000003810380010105C00102000040003C0FE7F0240E0F000C00000,
    pm.ram00_07.INIT_3C = 256'h383838387C7C7C7C8E387C7C7C7C7C7C5C383810000008001400005C0000007C,
    pm.ram00_07.INIT_3D = 256'h38383838383838386E383C3C3C3C3C3C20583810383878383800383838387044,
    pm.ram00_07.INIT_3E = 256'h000000000000000000000FF000F0000040043804383880383800383838383844,
    pm.ram00_07.INIT_3F = 256'h0000200000000000000000000000000000000000000000000000000000000000;
defparam
    pm.ram08_0F.INIT_00 = 256'h0000000000000000000000000000000000000000002000000000000000000000,
    pm.ram08_0F.INIT_01 = 256'h0000000070000000003C00000000000000000000000000000000000000000006,
    pm.ram08_0F.INIT_02 = 256'h00FF0000000000000201080420108040005500000000003C0000000000006006,
    pm.ram08_0F.INIT_03 = 256'h00000000000000000000000000000000200004000180FFFF0180E0F000C00000,
    pm.ram08_0F.INIT_04 = 256'h0000000000000000006044444444444404000838000010000000004000000000,
    pm.ram08_0F.INIT_05 = 256'h0000000000000000006000000000000000800000000000000000000000000000,
    pm.ram08_0F.INIT_06 = 256'h401A40606203401A405A4050401A405D40380038000000000000000000000000,
    pm.ram08_0F.INIT_07 = 256'h401A405A62034050401A40634058401A405D720F4056401A406362034066720F,
    pm.ram08_0F.INIT_08 = 256'h612340636203401A40638001403E4477401B4471401B4468720F6600FFFF6203,
    pm.ram08_0F.INIT_09 = 256'h401A405A8001448444844484448444844484448444846103612340638000710F,
    pm.ram08_0F.INIT_0A = 256'h44A444A40491449144914491449144914491449144914491710F6123405A6203,
    pm.ram08_0F.INIT_0B = 256'h405D6203401A405D800161036123405A800044AE04A444A444A444A444A444A4,
    pm.ram08_0F.INIT_0C = 256'h405A800004B644C244C244C204B644B644B644B644B644B644B644B6710F6123,
    pm.ram08_0F.INIT_0D = 256'h89C20000700C89BC720F804044D7700CBF0004CA61036123405D800061036123,
    pm.ram08_0F.INIT_0E = 256'h801840048000401A44DF6103612344DC400F804F40048000401A44DC0000700C,
    pm.ram08_0F.INIT_0F = 256'h04E2404444DF6600800004E26103612344DC6103612344DF710F612344DF400F,
    pm.ram08_0F.INIT_10 = 256'h4058401A44DF04E2404444DC800104E2404444DC6600800004E2404444DF8001,
    pm.ram08_0F.INIT_11 = 256'h8050403E61806600401B608160810000700C8A30720F6600FFFF6203401A44DC,
    pm.ram08_0F.INIT_12 = 256'h650366008000401A4516610345194519451945194519451945194519450D720F,
    pm.ram08_0F.INIT_13 = 256'h60816203401A453880010000700C8A74700C45212537401A4516710F61234516,
    pm.ram08_0F.INIT_14 = 256'h0000700C8A9E710F61234538800045216103710F61234538254765036600BFFF,
    pm.ram08_0F.INIT_15 = 256'h002300210032001C0046003E003D0036002E00250026001E00160045700C8AA4,
    pm.ram08_0F.INIT_16 = 256'h004200410039003800370036003500340033003200310030700C8AC8002B0024,
    pm.ram08_0F.INIT_17 = 256'h000B006A0C0000BF000B006A130000CF000B006A700C8AEC0046004500440043,
    pm.ram08_0F.INIT_18 = 256'h000B0070140000EF000B00701200000F000B006D0C0000BF000B006D060000BF,
    pm.ram08_0F.INIT_19 = 256'h000B0071060000BF000B00711200000F000B00704400008F000B0070110000EF,
    pm.ram08_0F.INIT_1A = 256'h000B0071060000DF000B0071180000EF000B0071190000CF000B00710D00005F,
    pm.ram08_0F.INIT_1B = 256'h000B00730D00005F000B0073060000FF000B00710D00005F000B0071130000CF,
    pm.ram08_0F.INIT_1C = 256'h000B0077110000CF000B00771300000F000B00740C0000BF000B0074060000FF,
    pm.ram08_0F.INIT_1D = 256'h000B007A1200004F000B007A440000AF000B00794500003F000B00771700002F,
    pm.ram08_0F.INIT_1E = 256'h000B007B440000AF000B007A4500003F000B007A1700000F000B007A1200002F,
    pm.ram08_0F.INIT_1F = 256'h000B007C460000FF000B007B4500003F000B007B1700002F000B007B110000CF,
    pm.ram08_0F.INIT_20 = 256'h000B007D4600004F000B007D4500003F000B007D1200004F000B007D440000AF,
    pm.ram08_0F.INIT_21 = 256'h000B007E4600004F000B007E450000FF000B007E1200004F000B007E440000AF,
    pm.ram08_0F.INIT_22 = 256'h000B0080450000FF000B00804500003F000B00801200000F000B0080430000FF,
    pm.ram08_0F.INIT_23 = 256'h000B008B0F00009F000B008A0F00007F000B008A440000AF000B008A0F00009F,
    pm.ram08_0F.INIT_24 = 256'h000B008C1200002F000B008C1700002F000B008C1300000F000B008C1200002F,
    pm.ram08_0F.INIT_25 = 256'h000B008D110000EF000B008D140000EF000B008D1B0000FF000B008D120000AF,
    pm.ram08_0F.INIT_26 = 256'h000B008E1700000F000B008E0F00009F000B008E1200002F000B008E0F00007F,
    pm.ram08_0F.INIT_27 = 256'h000B00911200000F000B00910F00007F000B0090110000EF000B008E0F00009F,
    pm.ram08_0F.INIT_28 = 256'h000B0093120000CF000B00930F00007F000B00921700002F000B00921300000F,
    pm.ram08_0F.INIT_29 = 256'h000B00970F00009F000B0097470000DF000B00971200000F000B00944500003F,
    pm.ram08_0F.INIT_2A = 256'h000B00971700000F000B00971200002F000B00970F00007F000B0097440000AF,
    pm.ram08_0F.INIT_2B = 256'h000B009A0F00007F000B009A440000AF000B009A0F00009F000B00974500003F,
    pm.ram08_0F.INIT_2C = 256'h000B009B120000EF000B009B120000AF000B009B120000AF000B009A120000AF,
    pm.ram08_0F.INIT_2D = 256'h000B009C110000CF000B009B1300006F000B009B120000AF000B009B140000EF,
    pm.ram08_0F.INIT_2E = 256'h000E002D5000001F000E002D120000CF000C00534A00001F000C00530E00005F,
    pm.ram08_0F.INIT_2F = 256'h000E0032370000CF000E00324400005F000E002E5000004F000E002E120000CF,
    pm.ram08_0F.INIT_30 = 256'h000E00341200000F000E00331300000F000E00333500009F000E0032180000AF,
    pm.ram08_0F.INIT_31 = 256'h000E00351200002F000E00343A0000EF000E00341200000F000E00343900001F,
    pm.ram08_0F.INIT_32 = 256'h000E00350D00005F000E00351200002F000E00354A0000EF000E00351700000F,
    pm.ram08_0F.INIT_33 = 256'h000E003B1200000F000E003A1300000F000E003A3500009F000E00394A00005F,
    pm.ram08_0F.INIT_34 = 256'h000E003C3A0000EF000E003C1200000F000E003B3500009F000E003B180000AF,
    pm.ram08_0F.INIT_35 = 256'h000E003D3500009F000E003D180000AF000E003D180000AF000E003D1200000F,
    pm.ram08_0F.INIT_36 = 256'h000E003E4B00000F000E003E1700000F000E003E120000AF000E003D0C0000BF,
    pm.ram08_0F.INIT_37 = 256'h000E004351000075000E00435100000A000E003F0D00005F000E003F1200002F,
    pm.ram08_0F.INIT_38 = 256'h000F000D1300004F000F000D1600008F000F000D1200000F000F000D4D0000AF,
    pm.ram08_0F.INIT_39 = 256'h000F00101300004F000F00101600008F000F00101200000F000F00104D0000DF,
    pm.ram08_0F.INIT_3A = 256'h001000371200000F001000251300006F000F0012110000EF000F00124C0000CF,
    pm.ram08_0F.INIT_3B = 256'h001000371800002F001000371200002F001000371300006F001000371300004F,
    pm.ram08_0F.INIT_3C = 256'h001000380F0000BF001000381100007F001000381C00001F001000371300006F,
    pm.ram08_0F.INIT_3D = 256'h001000394E00009F00100039120000CF001000390F00007F001000382C0000BF,
    pm.ram08_0F.INIT_3E = 256'h0010003C1300004F001000391300004F00100039160000CF001000391200000F,
    pm.ram08_0F.INIT_3F = 256'h0010003C2C0000BF0010003C0F0000BF0010003C1100007F0010003C1C00001F;
defparam
    pm.ram10_17.INIT_00 = 256'h0010003D1200000F0010003D4E00009F0010003D120000CF0010003D0F00007F,
    pm.ram10_17.INIT_01 = 256'h0010003F1600006F0010003F4E0000CF0010003D1300004F0010003D160000CF,
    pm.ram10_17.INIT_02 = 256'h001000422C0000BF001000420F0000BF001000421100007F0010003F1300004F,
    pm.ram10_17.INIT_03 = 256'h001000421300004F001000421600006F001000424C00007F001000420F00007F,
    pm.ram10_17.INIT_04 = 256'h001000450F00007F001000452C0000BF001000450F0000BF001000451100007F,
    pm.ram10_17.INIT_05 = 256'h001000452C0000BF001000450F0000BF001000451100007F00100045120000CF,
    pm.ram10_17.INIT_06 = 256'h001000451600006F001000454C0000EF001000451200002F001000450F00007F,
    pm.ram10_17.INIT_07 = 256'h001000531200000F001000534F00002F00100053120000CF001000451300004F,
    pm.ram10_17.INIT_08 = 256'h001000531300004F00100053160000CF001000531200002F00100053150000AF,
    pm.ram10_17.INIT_09 = 256'h001000561300004F00100056160000CF001000564E0000FF00100056120000CF,
    pm.ram10_17.INIT_0A = 256'h0010006D1100007F001000591300004F00100059160000CF001000594D00001F,
    pm.ram10_17.INIT_0B = 256'h0010006D5700004F0010006D0F00007F0010006D500000BF0010006D0F0000BF,
    pm.ram10_17.INIT_0C = 256'h0010006D1600006F0010006D120000AF0010006D0C0000BF0010006D130000CF,
    pm.ram10_17.INIT_0D = 256'h00100074160000CF001000741200004F001000744F0000EF0010006D1300004F,
    pm.ram10_17.INIT_0E = 256'h00100077020000CF001000771B0000DF001000771200002F001000741300004F,
    pm.ram10_17.INIT_0F = 256'h001000781300004F00100078160000CF001000784F0000EF001000781200002F,
    pm.ram10_17.INIT_10 = 256'h0010007C1200002F0010007B020000CF0010007B1B0000DF0010007B1200002F,
    pm.ram10_17.INIT_11 = 256'h0010007F1100007F0010007C1300004F0010007C1600006F0010007C4D00004F,
    pm.ram10_17.INIT_12 = 256'h0010007F1200000F0010007F0F0000BF0010007F2C0000BF0010007F0F0000BF,
    pm.ram10_17.INIT_13 = 256'h0010007F1200002F0010007F0D00001F0010007F0F00007F0010007F5000007F,
    pm.ram10_17.INIT_14 = 256'h001000A05700006F001000A01200000F0010007F1300004F0010007F160000CF,
    pm.ram10_17.INIT_15 = 256'h001000A01B0000DF001000A0110000EF001000A00F00009F001000A01300000F,
    pm.ram10_17.INIT_16 = 256'h001000A11200002F001000A0110000EF001000A0020000CF001000A00F00007F,
    pm.ram10_17.INIT_17 = 256'h93020000700C92FC0000700C92F60000700C92F01200004F001000A10F00009F,
    pm.ram10_17.INIT_18 = 256'h66008000618062038001403E618180206180299260810000700C93080000700C,
    pm.ram10_17.INIT_19 = 256'h710F612344DF80006103612344DC8000498587D0401A4060710F610309856203,
    pm.ram10_17.INIT_1A = 256'h450949A4003E62036203401A44DC4050401A44DF401A4060710F612340604574,
    pm.ram10_17.INIT_1B = 256'h62038001618062036600800049AE401B618129C26081710F6123497666008000,
    pm.ram10_17.INIT_1C = 256'h09D86303800F09AE802B09AE802005006103612344DC8000710F610309B56180,
    pm.ram10_17.INIT_1D = 256'h8004608109AE401B62036103801093A045464344414238393637343532333031,
    pm.ram10_17.INIT_1E = 256'h49E949E9720F800249E3401A608109C949DE49DE69038008608109CD49CD6903,
    pm.ram10_17.INIT_1F = 256'h49F649F649F649F649F6720F800149AE401B608109E949E949E949E949E949E9,
    pm.ram10_17.INIT_20 = 256'h941A20202D2D0A0F49EE09F649F649F649F649F649F649F649F649F649F649F6,
    pm.ram10_17.INIT_21 = 256'h6E20656550726C20726573744B650A21710F49C449FB62036600800F49B58003,
    pm.ram10_17.INIT_22 = 256'h0A0BBF0049B58007944E202430202030442B0A2B09C449C449B5801094323141,
    pm.ram10_17.INIT_23 = 256'h9476202730202032442B0A3F0A0BBF1049B580079462208F30202031442B0A35,
    pm.ram10_17.INIT_24 = 256'h4A304A260A0BBF3049B58007948A206F30202033442B0A490A0BBF2049B58007,
    pm.ram10_17.INIT_25 = 256'h2031522B0A620A0BBF3F49B5800794A8201230202030522B0A5809C44A444A3A,
    pm.ram10_17.INIT_26 = 256'hBF6049B5800794D0201230202032522B0A6C0A0BBF5049B5800794BC20003020,
    pm.ram10_17.INIT_27 = 256'h09C44A714A674A5D4A530A0BBF7049B5800794E4200030202033522B0A760A0B,
    pm.ram10_17.INIT_28 = 256'h401A4A80608149C949C949DE608149B58003950820004D2B0A860000700C9504,
    pm.ram10_17.INIT_29 = 256'h4A83800049C449E3401A4A8049B58003952A204E4D3D0A97720F80104A0B6203,
    pm.ram10_17.INIT_2A = 256'h474F0AB04A944A7B4A4E4A18499409C461034A834A834A834A834A834A834A83,
    pm.ram10_17.INIT_2B = 256'h6103610349AE4AB4001A620345626203800162036600455009C449B58002955E,
    pm.ram10_17.INIT_2C = 256'h4AC1710F6B8D6B8D610361036B8D6B8D4ABC700C2AC76503401A61816181710F,
    pm.ram10_17.INIT_2D = 256'h4ACF4ACF4ACF4ACF4ACF4ACF4ACF4ACF4ACF4ACF4ACF4ACF4ACF4ACF720F8002,
    pm.ram10_17.INIT_2E = 256'h710F61036B8D44FB700C2AEC650381756081710F61034AD2455060810ACF4ACF,
    pm.ram10_17.INIT_2F = 256'h6B8D4504700C2AFE6503816B6081710F61036B8D4500700C2AF5650381726081,
    pm.ram10_17.INIT_30 = 256'h720F401A497C401A4982710F61036B8D4509700C2B07650381746081710F6103,
    pm.ram10_17.INIT_31 = 256'h710F6B8D700C2B1E63036600FFFF62038001620366008050401A4982001B4B0B,
    pm.ram10_17.INIT_32 = 256'h0B294044498280012B304B204B12730F6600FFFF620380016203660080214B10,
    pm.ram10_17.INIT_33 = 256'h6203660061814B0B4B314B0B4B290B31404449828001700C2B354B204B12700C,
    pm.ram10_17.INIT_34 = 256'h2B5163036600FFFF620366008009608162036600802F0000700C9688720F8001,
    pm.ram10_17.INIT_35 = 256'h6081710F61234B4264036D038004401A4B424B45401B6181720F66008006700C,
    pm.ram10_17.INIT_36 = 256'h610361234B428000710F61030B5F61806203800161806203660080004B542B6A,
    pm.ram10_17.INIT_37 = 256'h4B744B744B744B744B744B74720F80026103612361814B6C001A4B424B5F4B39,
    pm.ram10_17.INIT_38 = 256'h610361234A804B6C0B7A620344D94B6C0B7A620344D74B6C0AA961034B744B74,
    pm.ram10_17.INIT_39 = 256'hBF786147401ABF7A6147401ABF7C6147401ABF7E0B7A6203401A4A804B6C0AA9,
    pm.ram10_17.INIT_3A = 256'h401ABF6E6147401ABF706147401ABF726147401ABF746147401ABF766147401A,
    pm.ram10_17.INIT_3B = 256'h6147401ABF646147401ABF666147401ABF686147401ABF6A6147401ABF6C6147,
    pm.ram10_17.INIT_3C = 256'hBF586147401ABF5A6147401ABF5C6147401ABF5E6147401ABF606147401ABF62,
    pm.ram10_17.INIT_3D = 256'h401ABF4E6147401ABF506147401ABF526147401ABF546147401ABF566147401A,
    pm.ram10_17.INIT_3E = 256'h6147401ABF446147401ABF466147401ABF486147401ABF4A6147401ABF4C6147,
    pm.ram10_17.INIT_3F = 256'h401ABF36401ABF38401ABF3A401ABF3C401ABF3E6147401ABF3F6147401ABF42;
defparam
    pm.ram18_1F.INIT_00 = 256'h401ABF26401ABF28401ABF2A401ABF2C401ABF2E401ABF30401ABF32401ABF34,
    pm.ram18_1F.INIT_01 = 256'h401ABF16401ABF18401ABF1A401ABF1C401ABF1E401ABF20401ABF22401ABF24,
    pm.ram18_1F.INIT_02 = 256'h401ABF06401ABF08401ABF0A401ABF0C401ABF0E401ABF10401ABF12401ABF14,
    pm.ram18_1F.INIT_03 = 256'h442B700C987E0B960B910B8C0B880B84700C9870001ABF00401ABF02401ABF04,
    pm.ram18_1F.INIT_04 = 256'h6181001A62034C3662038001620366004C3D0AA9700C988C474F4D2B4D3D522B,
    pm.ram18_1F.INIT_05 = 256'h4C4F4C4F4C3D710F61036B8D6B8D4C4761036180720F80022C566503401A6181,
    pm.ram18_1F.INIT_06 = 256'h4B39710F6B8D700C2C6D6081001A4C4461034C5D401A6103700C4C4F4C4F4C4F,
    pm.ram18_1F.INIT_07 = 256'h6123497F805061036123497C6203401A40604050401A44DF700C61474C644C6A,
    pm.ram18_1F.INIT_08 = 256'h4AE7710F61036B8D4C74700C2C8B6503805A60810C6F61036123498280006103,
    pm.ram18_1F.INIT_09 = 256'h454D8100700C2C9E650380E0608105214C8F4533710F4AE24C864B024AF94AF0,
    pm.ram18_1F.INIT_0A = 256'h454D6600FFFF700C2CAD650380F06081710F61036B8D61036123454D6403401A,
    pm.ram18_1F.INIT_0B = 256'h454D80004C966403401A454D4CA84C99710F61036B8D61036123454D6403401A,
    pm.ram18_1F.INIT_0C = 256'h660080018300730F80FF401A66008001730F6600FFFF401A66008001710F6123,
    pm.ram18_1F.INIT_0D = 256'h49768000452144CE45332CE2401A4976700C4CCD4CB84CC82CD74CC2710F6123,
    pm.ram18_1F.INIT_0E = 256'h800061036123454D8000700C0CE32CEA401A49794CD2453B4CD8700C61036123,
    pm.ram18_1F.INIT_0F = 256'hBF0661036123BF0461036123BF0261036123BF0005334CE36103612349796600,
    pm.ram18_1F.INIT_10 = 256'h6123BF1061036123BF0E61036123BF0C61036123BF0A61036123BF0861036123,
    pm.ram18_1F.INIT_11 = 256'h61036123BF1A61036123BF1861036123BF1661036123BF1461036123BF126103,
    pm.ram18_1F.INIT_12 = 256'hBF2661036123BF2461036123BF2261036123BF2061036123BF1E61036123BF1C,
    pm.ram18_1F.INIT_13 = 256'h6123BF3061036123BF2E61036123BF2C61036123BF2A61036123BF2861036123,
    pm.ram18_1F.INIT_14 = 256'h61036123BF3A61036123BF3861036123BF3661036123BF3461036123BF326103,
    pm.ram18_1F.INIT_15 = 256'hBF446B8D61036123BF426B8D61036123BF3F6B8D61036123BF3E61036123BF3C,
    pm.ram18_1F.INIT_16 = 256'hBF4C6B8D61036123BF4A6B8D61036123BF486B8D61036123BF466B8D61036123,
    pm.ram18_1F.INIT_17 = 256'hBF546B8D61036123BF526B8D61036123BF506B8D61036123BF4E6B8D61036123,
    pm.ram18_1F.INIT_18 = 256'hBF5C6B8D61036123BF5A6B8D61036123BF586B8D61036123BF566B8D61036123,
    pm.ram18_1F.INIT_19 = 256'hBF646B8D61036123BF626B8D61036123BF606B8D61036123BF5E6B8D61036123,
    pm.ram18_1F.INIT_1A = 256'hBF6C6B8D61036123BF6A6B8D61036123BF686B8D61036123BF666B8D61036123,
    pm.ram18_1F.INIT_1B = 256'hBF746B8D61036123BF726B8D61036123BF706B8D61036123BF6E6B8D61036123,
    pm.ram18_1F.INIT_1C = 256'hBF7C6B8D61036123BF7A6B8D61036123BF786B8D61036123BF766B8D61036123,
    pm.ram18_1F.INIT_1D = 256'h0014002E1200000F0014700C9BB60CEB4AA949A061036123BF7E6B8D61036123,
    pm.ram18_1F.INIT_1E = 256'h0014002F1200000F0014002E020000CF0014002E6A0000310014002E140000EF,
    pm.ram18_1F.INIT_1F = 256'h001400301200000F0014002F020000CF0014002F6A0000AB0014002F140000EF,
    pm.ram18_1F.INIT_20 = 256'h001400316A0000D000140030020000CF001400306A00007900140030140000EF,
    pm.ram18_1F.INIT_21 = 256'h00140035160000AF00140035160000CF001400351200000F001400341200002F,
    pm.ram18_1F.INIT_22 = 256'h001400396B0000E9001400371B0000DF001400366B000038001400362500002F,
    pm.ram18_1F.INIT_23 = 256'h0014004E0C0000BF0014004E070000EF0014003B0C0000BF0014003B0600007F,
    pm.ram18_1F.INIT_24 = 256'h001400510800002F001400511500008F001400511700000F001400516C00008F,
    pm.ram18_1F.INIT_25 = 256'h001400530600005F001400511300004F001400511600008F001400510C0000BF,
    pm.ram18_1F.INIT_26 = 256'h001400580800004F001400586D00001F001400556C0000EF001400530E00005F,
    pm.ram18_1F.INIT_27 = 256'h001400730E0000DF001400730800004F001400582A00007F001400580C0000BF,
    pm.ram18_1F.INIT_28 = 256'h001400732600006F00140073090000AF001400730C0000BF001400730600007F,
    pm.ram18_1F.INIT_29 = 256'h001400760800004F001400736100002F001400730D00005F001400730600005F,
    pm.ram18_1F.INIT_2A = 256'h001400766D00009F001400760C0000BF001400760800002F001400760E0000DF,
    pm.ram18_1F.INIT_2B = 256'h001400796E00002F001400791700000F001400796C00008F001400766D00006F,
    pm.ram18_1F.INIT_2C = 256'h0014007C6C00008F0014007B0E0000DF0014007B080000AF0014007B300000EF,
    pm.ram18_1F.INIT_2D = 256'h0015002470000038001500246F00005F0014007C6D0000CF0014007C6E00007F,
    pm.ram18_1F.INIT_2E = 256'h001500250D00005F0015002570000038001500256F00007F001500240D00005F,
    pm.ram18_1F.INIT_2F = 256'h0015002A0D00003F0015002A130000CF0015002A6F0000AA0015002A0D00003F,
    pm.ram18_1F.INIT_30 = 256'h001500531600008F001500534E00006F001500536F0000AA001500536F00003F,
    pm.ram18_1F.INIT_31 = 256'h001500546F0000F1001500546F0000AA001500530D00005F001500536F00009F,
    pm.ram18_1F.INIT_32 = 256'h001500550E00005F001500551200000F00150055720000A7001500542900002F,
    pm.ram18_1F.INIT_33 = 256'h001500550C0000BF00150055130000CF00150055190000CF001500556F0000F1,
    pm.ram18_1F.INIT_34 = 256'h00150056190000CF001500566F0000F1001500551300006F001500551300004F,
    pm.ram18_1F.INIT_35 = 256'h00150056110000EF00150056130000CF001500560D00005F00150056130000CF,
    pm.ram18_1F.INIT_36 = 256'h00150059110000EF001500594E00006F001500596F0000AA001500596F00003F,
    pm.ram18_1F.INIT_37 = 256'h0015005E110000EF0015005E4E00006F0015005E6F0000F10015005E6F00003F,
    pm.ram18_1F.INIT_38 = 256'h0015006C730000C90015006C0C0000BF0015006C6F00009F0015006C2300005F,
    pm.ram18_1F.INIT_39 = 256'h0015006D4C00002F0015006D0C0000BF0015006D7400003F0015006C260000AF,
    pm.ram18_1F.INIT_3A = 256'h00150070110000EF001500704E0000FF00150070120000CF001500706F00007F,
    pm.ram18_1F.INIT_3B = 256'h001500864F00005F0015008675000005001500727400005F001500707400005F,
    pm.ram18_1F.INIT_3C = 256'h001500894F00002F00150089740000FA001500896F00003F001500861400002F,
    pm.ram18_1F.INIT_3D = 256'h0015008C70000038001500890D00003F00150089740000FA00150089110000EF,
    pm.ram18_1F.INIT_3E = 256'h0015008C110000EF0015008C4E0000FF0015008C120000CF0015008C0C0000BF,
    pm.ram18_1F.INIT_3F = 256'h0015008F0C0000BF0015008F700000380015008F0D00009F0015008F740000FA;
defparam
    pm.ram20_27.INIT_00 = 256'h001500911100007F0015008F110000EF0015008F4E0000FF0015008F740000FA,
    pm.ram20_27.INIT_01 = 256'h00150092110000EF001500924E00006F001500920F0000BF001500926F00003F,
    pm.ram20_27.INIT_02 = 256'h001500A47500008A001500931A00009F001500930C0000BF001500930F00007F,
    pm.ram20_27.INIT_03 = 256'h001500A80F00009F001500A80C0000BF001500A80600009F001500A62200009F,
    pm.ram20_27.INIT_04 = 256'h001500A96700006F001500A91700000F001500A87600000C001500A8610000FF,
    pm.ram20_27.INIT_05 = 256'h001500A90600009F001500A90F00007F001500A96700006F001500A91700000F,
    pm.ram20_27.INIT_06 = 256'h001500AC1600002F001500AC1200000F001500AC2400002F001500A90D00005F,
    pm.ram20_27.INIT_07 = 256'h001500AC130000CF001500AC3C00004F001500AC1200002F001500AC1400000F,
    pm.ram20_27.INIT_08 = 256'h001500B07600000C001500AD1700002F001500AD1300000F001500AD110000EF,
    pm.ram20_27.INIT_09 = 256'h001500B1140000EF001500B12400002F001500B0140000EF001500B02400002F,
    pm.ram20_27.INIT_0A = 256'h001500B11200002F001500B17600009A001500B17600009A001500B11B0000DF,
    pm.ram20_27.INIT_0B = 256'h001500B4110000CF001500B4750000BF001500B4110000CF001500B477000036,
    pm.ram20_27.INIT_0C = 256'h001500B5750000F9001500B51700000F001500B4250000AF001500B41700002F,
    pm.ram20_27.INIT_0D = 256'h001500BF0F00009F001500BF0C0000BF001500BF0600009F001500B5250000AF,
    pm.ram20_27.INIT_0E = 256'h001500BF78000021001500BF150000CF001500BF150000AF001500BF610000FF,
    pm.ram20_27.INIT_0F = 256'h001500C01300000F001500BF7600000C001500BF0D00003F001500BF130000CF,
    pm.ram20_27.INIT_10 = 256'h001500C0140000CF001500C0220000DF001500C06500008F001500C01200000F,
    pm.ram20_27.INIT_11 = 256'h001500CA1200004F001500C10D00005F001500C10600009F001500C10F00007F,
    pm.ram20_27.INIT_12 = 256'h001500CA4F00002F001500CA1200004F001500CA6F00003F001500CA1200002F,
    pm.ram20_27.INIT_13 = 256'h001500CB1700000F001500CB140000EF001500CB0D00003F001500CB1200000F,
    pm.ram20_27.INIT_14 = 256'h001500CD1200002F001500CC740000EF001500CC1600008F001500CC190000CF,
    pm.ram20_27.INIT_15 = 256'h001500D04F00002F001500D0740000FA001500D06F00003F001500CD1400000F,
    pm.ram20_27.INIT_16 = 256'h001500D00D00003F001500D0740000FA001500D0740000EF001500D01600008F,
    pm.ram20_27.INIT_17 = 256'h001500E47500008A001500E31300002F001500E21300002F001500E11300002F,
    pm.ram20_27.INIT_18 = 256'h001500E8770000C0001500E7750000F9001500E675000067001500E575000067,
    pm.ram20_27.INIT_19 = 256'h001500EC75000039001500EB75000014001500EA75000039001500E97800002D,
    pm.ram20_27.INIT_1A = 256'h001500F07600002C001500EF1B0000DF001500EE75000039001500ED75000014,
    pm.ram20_27.INIT_1B = 256'h001500FA1300002F001500F36C00004F001500F2750000BF001500F177000036,
    pm.ram20_27.INIT_1C = 256'h001500FE75000067001500FD7500008A001500FC1300002F001500FB1300002F,
    pm.ram20_27.INIT_1D = 256'h62038001403E6181618100011300002F01150000750000F9001500FF75000067,
    pm.ram20_27.INIT_1E = 256'h51DB51DB51DB51DB51DB51DB51DB51DB51DB51DB51DB51DB718C620380016180,
    pm.ram20_27.INIT_1F = 256'h51F451F451F451F451F451F451F4720F8001403E6181802011DB51DB51DB51DB,
    pm.ram20_27.INIT_20 = 256'h520D120951E411F951F951F951F911F451F451F451F451F451F451F451F451F4,
    pm.ram20_27.INIT_21 = 256'h802E120D520D520D520D520D520D520D520D520D520D520D520D520D520D520D,
    pm.ram20_27.INIT_22 = 256'h52245224121F521F521F521F521F521F521F521F521F521F720F8001403E6181,
    pm.ram20_27.INIT_23 = 256'h8000122E522E522E522E522E522E522E522E522E122452245224522452245224,
    pm.ram20_27.INIT_24 = 256'h4DD9523F1245610361236600FEFF6600401A6600FEFF710F61035236520F4DD9,
    pm.ram20_27.INIT_25 = 256'h12574CF61257610361236600F777660080001245601044CE6010610361234060,
    pm.ram20_27.INIT_26 = 256'h001600226D00003F0016001F0E00007F0016001F0800004F0016001F130000CF,
    pm.ram20_27.INIT_27 = 256'h001600222A0000EF001600221B00002F001600220F00009F001600221200004F,
    pm.ram20_27.INIT_28 = 256'h001600220800004F001600221400000F001600220F00007F00160022110000EF,
    pm.ram20_27.INIT_29 = 256'h001600230600007F00160023110000EF001600236D00003F001600220E00007F,
    pm.ram20_27.INIT_2A = 256'h001600230D00005F00160023080000CF001600231400000F001600230C0000BF,
    pm.ram20_27.INIT_2B = 256'h00160023180000AF00160023080000CF001600231200000F001600237B0000AF,
    pm.ram20_27.INIT_2C = 256'h001600245D00006F001600240D00009F001600245D00006F001600230D00005F,
    pm.ram20_27.INIT_2D = 256'h001600276D00003F001600245D00006F001600242900002F001600242900000F,
    pm.ram20_27.INIT_2E = 256'h001600272A0000EF001600270900000F001600270F00009F001600271200004F,
    pm.ram20_27.INIT_2F = 256'h001600270800004F001600271400000F001600270F00007F00160027110000EF,
    pm.ram20_27.INIT_30 = 256'h0017007F0000003F001600277B0000AF001600270900000F001600270E00007F,
    pm.ram20_27.INIT_31 = 256'h0017007F7E00004F0017007F0F00009F0017007F1200002F0017007F0F00001F,
    pm.ram20_27.INIT_32 = 256'h0017008B0C0000BF0017008B0A0000DF0017007F130000CF0017007F0F00007F,
    pm.ram20_27.INIT_33 = 256'h0017008B1300006F0017008B1800004F0017008B0C0000BF0017008B0A0000FF,
    pm.ram20_27.INIT_34 = 256'h0017008B0E00002F0017008B0C0000BF0017008B7E0000EF0017008B1200002F,
    pm.ram20_27.INIT_35 = 256'h0017008E1200000F0017008E130000CF0017008B0E00007F0017008B7E0000EF,
    pm.ram20_27.INIT_36 = 256'h0017008F3500009F0017008F7E0000FE0017008E0E00002F0017008E7E0000EF,
    pm.ram20_27.INIT_37 = 256'h0017008F0F00009F0017008F0F00001F0017008F1200000F0017008F1300000F,
    pm.ram20_27.INIT_38 = 256'h001700902900002F001700900F0000BF001700900C0000BF001700907E0000EF,
    pm.ram20_27.INIT_39 = 256'h001700912A00001F00170091180000AF001700910C0000BF001700911200000F,
    pm.ram20_27.INIT_3A = 256'h001700927E0000FE001700920E00007F001700927E0000EF001700920F00007F,
    pm.ram20_27.INIT_3B = 256'h001700AD1200006F001700AC1200004F001700947F000009001700920D00005F,
    pm.ram20_27.INIT_3C = 256'h001700AD7D0000DF001700AD7E00009F001700AD120000AF001700AD1200006F,
    pm.ram20_27.INIT_3D = 256'h001700AE020000CF001700AD8000004F001700AD1200004F001700AD1200000F,
    pm.ram20_27.INIT_3E = 256'h001700B20C0000BF001700B2060000BF001700B2060000DF001700AF4100007F,
    pm.ram20_27.INIT_3F = 256'h001700B21200002F001700B2130000CF001700B21200004F001700B2180000EF;
defparam
    pm.ram28_2F.INIT_00 = 256'h001700B38000007F001700B30C0000BF001700B3190000CF001700B31B0000FF,
    pm.ram28_2F.INIT_01 = 256'h001700B3020000CF001700B3190000AF001700B31C00007F001700B31300000F,
    pm.ram28_2F.INIT_02 = 256'h001700B72900000F001700B71200000F001700B41B0000DF001700B41800006F,
    pm.ram28_2F.INIT_03 = 256'h001700B8120000AF001700B81200000F001700B88100000F001700B71200000F,
    pm.ram28_2F.INIT_04 = 256'h001700BC0900000F001700B91B0000DF001700B8020000CF001700B8110000EF,
    pm.ram28_2F.INIT_05 = 256'h001700BE110000CF001700BE8200003F001700BC810000BF001700BC7C00005F,
    pm.ram28_2F.INIT_06 = 256'h001800270C0000BF001800270A00006F001700BF160000AF001700BF8200006F,
    pm.ram28_2F.INIT_07 = 256'h00180027110000EF00180027020000CF001800271700002F001800271200000F,
    pm.ram28_2F.INIT_08 = 256'h0018002A1300004F0018002A0D00003F0018002A820000CB001800275D00006F,
    pm.ram28_2F.INIT_09 = 256'h0018002C820000F60018002A0D00009F0018002A820000CB0018002A1300006F,
    pm.ram28_2F.INIT_0A = 256'h00180030390000DF001800302300005F0018002E820000F60018002D820000F6,
    pm.ram28_2F.INIT_0B = 256'h001800330C00006F00180033830000BD00180030220000DF001800302900000F,
    pm.ram28_2F.INIT_0C = 256'h0018003A4100009F001800393100001F00180036830000BD001800330E0000FF,
    pm.ram28_2F.INIT_0D = 256'h0018003C0C00007A0018003B3100001F0018003A830000DC0018003A8000007F,
    pm.ram28_2F.INIT_0E = 256'h0018003D0E0000BF0018003D0C00007A0018003C1600008F0018003C0C0000BF,
    pm.ram28_2F.INIT_0F = 256'h0018003F0C00007A0018003E8400000D0018003E8000007F0018003E4100009F,
    pm.ram28_2F.INIT_10 = 256'h0018004D0A0000DF0018004D6C0000AF00180043300000EF0018003F0E0000DF,
    pm.ram28_2F.INIT_11 = 256'h0018004D0C0000BF0018004D0A0000FF0018004D150000CF0018004D0C0000BF,
    pm.ram28_2F.INIT_12 = 256'h001800511200000F001800517E00009F0018004D1300006F0018004D1800004F,
    pm.ram28_2F.INIT_13 = 256'h001800510D00005F00180051130000CF00180051180000EF001800510A00006F,
    pm.ram28_2F.INIT_14 = 256'h001800525D00006F001800523600001F001800523500009F001800521200000F,
    pm.ram28_2F.INIT_15 = 256'h001800555D00006F00180052350000BF001800521200002F001800521400000F,
    pm.ram28_2F.INIT_16 = 256'h001800551200004F001800555D00006F001800550D00005F001800550A00006F,
    pm.ram28_2F.INIT_17 = 256'h0018006F1200004F001800552B0000EF001800555D00008F001800551700000F,
    pm.ram28_2F.INIT_18 = 256'h00180070120000CF0018006F840000350018006F3100005F0018006F1600008F,
    pm.ram28_2F.INIT_19 = 256'h001800702B0000EF001800700F0000BF001800701100007F00180070150000CF,
    pm.ram28_2F.INIT_1A = 256'h001800710D00003F001800710F0000BF00180071130000CF001800715D00006F,
    pm.ram28_2F.INIT_1B = 256'h001800711400000F001800711200002F001800711300004F00180071130000CF,
    pm.ram28_2F.INIT_1C = 256'h001800720F0000BF001800725E00001F001800728500002F001800715D00008F,
    pm.ram28_2F.INIT_1D = 256'h001800735E00008F001800728500009F00180072120000AF001800722900000F,
    pm.ram28_2F.INIT_1E = 256'h001800748600002F001800742900000F001800740F00007F001800735E00008F,
    pm.ram28_2F.INIT_1F = 256'h001800750A00006F001800755D00006F001800751700000F001800755D00006F,
    pm.ram28_2F.INIT_20 = 256'h001800780900000F001800755E00008F001800750E00002F00180075180000AF,
    pm.ram28_2F.INIT_21 = 256'h001800788600007F001800784600002F001800782900000F001800787C00005F,
    pm.ram28_2F.INIT_22 = 256'h0018007E2300001F0018007E2900000F0018007E1300000F0018007B8600007F,
    pm.ram28_2F.INIT_23 = 256'h001800860E0000DF001800860C00007A001800808800005F0018007E6100002F,
    pm.ram28_2F.INIT_24 = 256'h001900140C0000BF001900148900007F001800870E0000BF001800870C00007A,
    pm.ram28_2F.INIT_25 = 256'h001900150100004F001900140E00002F001900148900007F001900141200004F,
    pm.ram28_2F.INIT_26 = 256'h001900181200002F001900155E00001F001900155D00008F001900156000007F,
    pm.ram28_2F.INIT_27 = 256'h001900341200004F001900340E00007F00190034050000BF001900341200000F,
    pm.ram28_2F.INIT_28 = 256'h001900351200000F001900351400000F001900342F00006F001900340D00003F,
    pm.ram28_2F.INIT_29 = 256'h00190036140000CF001900351200000F001900351300006F001900351600002F,
    pm.ram28_2F.INIT_2A = 256'h001900360600009F001900361200000F001900361400000F001900361300004F,
    pm.ram28_2F.INIT_2B = 256'h001900370F00009F001900371200002F001900361600002F001900360C0000BF,
    pm.ram28_2F.INIT_2C = 256'h001900373C00004F001900370C0000BF001900370600009F001900371C00001F,
    pm.ram28_2F.INIT_2D = 256'h001900373C00000F001900370C0000BF001900370600009F001900371200002F,
    pm.ram28_2F.INIT_2E = 256'h001900380F00007F001900371700000F00190037120000AF001900371D00002F,
    pm.ram28_2F.INIT_2F = 256'h00190038020000CF001900381600008F001900381200000F001900381700002F,
    pm.ram28_2F.INIT_30 = 256'h0019003B110000EF0019003B8A00006F0019003B1700000F00190038110000EF,
    pm.ram28_2F.INIT_31 = 256'h0019003E0D00003F0019003E1200004F0019003E0D00005F0019003E050000BF,
    pm.ram28_2F.INIT_32 = 256'h0019003E0D00005F0019003E8A00004F0019003E1200000F0019003E140000EF,
    pm.ram28_2F.INIT_33 = 256'h0019003F1B0000DF0019003F140000AF0019003F1200000F0019003E2A00007F,
    pm.ram28_2F.INIT_34 = 256'h001900401200000F001900408A00006F0019003F1C00001F0019003F020000CF,
    pm.ram28_2F.INIT_35 = 256'h001900411600002F001900411200000F001900410D00003F001900411200004F,
    pm.ram28_2F.INIT_36 = 256'h001900422A00007F001900421300006F00190042140000EF001900421200002F,
    pm.ram28_2F.INIT_37 = 256'h001900431B0000DF001900431B0000DF001900420D00005F00190042050000BF,
    pm.ram28_2F.INIT_38 = 256'h001900440C0000BF001900448A00004F001900441B0000DF00190043020000CF,
    pm.ram28_2F.INIT_39 = 256'h00190045160000CF001900450C0000BF00190045050000BF001900441D00005F,
    pm.ram28_2F.INIT_3A = 256'h001900451700002F001900450D00005F001900458A00004F001900451200002F,
    pm.ram28_2F.INIT_3B = 256'h00190048110000EF00190048140000EF001900481200000F001900471200002F,
    pm.ram28_2F.INIT_3C = 256'h00190049140000EF001900491200000F00190048020000CF00190048610000CF,
    pm.ram28_2F.INIT_3D = 256'h0019004A1200000F00190049020000CF00190049610000FF00190049110000EF,
    pm.ram28_2F.INIT_3E = 256'h0019004A020000CF0019004A6200002F0019004A110000EF0019004A140000EF,
    pm.ram28_2F.INIT_3F = 256'h0019004B6200005F0019004B110000EF0019004B140000EF0019004B1200000F;
defparam
    pm.ram30_37.INIT_00 = 256'h0019004F0600009F0019004C1700002F0019004C110000EF0019004B020000CF,
    pm.ram30_37.INIT_01 = 256'h0019004F0D00003F0019004F1200004F0019004F0F00009F0019004F0C0000BF,
    pm.ram30_37.INIT_02 = 256'h0019004F0F00007F0019004F8C00002F0019004F2A00007F0019004F8E00002E,
    pm.ram30_37.INIT_03 = 256'h001A001E0900000F001A001B1600008F0019004F0D00005F0019004F0600009F,
    pm.ram30_37.INIT_04 = 256'h001A001E8F0000BF001A001E0D00003F001A001E1200000F001A001E7C00005F,
    pm.ram30_37.INIT_05 = 256'h001A00240900000F001A00218F0000EF001A001E8F0000BF001A001E810000BF,
    pm.ram30_37.INIT_06 = 256'h001A00248F0000BF001A00240D00003F001A00241200000F001A00247C00005F,
    pm.ram30_37.INIT_07 = 256'h001A0024160000CF001A00248F0000BF001A00241200000F001A0024810000BF,
    pm.ram30_37.INIT_08 = 256'h001A002E1A0000FF001A00286000007F001A00288F0000EF001A00266000007F,
    pm.ram30_37.INIT_09 = 256'h001A00351B0000DF001A0030900000EF001A002E3100005F001A002E160000CF,
    pm.ram30_37.INIT_0A = 256'h001A003A1200000F001A003A9100005F001A003A1B0000FF001A00379100002A,
    pm.ram30_37.INIT_0B = 256'h001A003B1B0000FF001A003A110000EF001A003A020000CF001A003A1C00007F,
    pm.ram30_37.INIT_0C = 256'h001A003E1200000F001A003B1C00007F001A003B1200000F001A003B8100000F,
    pm.ram30_37.INIT_0D = 256'h001A003F8F00002F001A003F1B0000FF001A003E110000EF001A003E020000EF,
    pm.ram30_37.INIT_0E = 256'h001A0040110000CF001A0040140000EF001A003F0300002F001A003F1200000F,
    pm.ram30_37.INIT_0F = 256'h001A00408A00001F001A00401C00007F001A0040890000AF001A0040110000CF,
    pm.ram30_37.INIT_10 = 256'h001A0052200000EF001A00522B0000EF001A0052920000BF001A0043910000FF,
    pm.ram30_37.INIT_11 = 256'h001A00560300004F001A00566000007F001A0056160000CF001A0053930000DF,
    pm.ram30_37.INIT_12 = 256'h001A0059020000CF001A00599400002A001A00591200000F001A00599100007F,
    pm.ram30_37.INIT_13 = 256'h001A005A020000CF001A005A0300004F001A005A1200000F001A005A9200009F,
    pm.ram30_37.INIT_14 = 256'h001A005E0300004F001A005E9100007F001A005B9400001F001A005A110000EF,
    pm.ram30_37.INIT_15 = 256'h001A00609400001F001A005F020000EF001A005F9200009F001A005E020000CF,
    pm.ram30_37.INIT_16 = 256'h001A00710900000F001A00701600008F001A00700C0000BF001A00700800008F,
    pm.ram30_37.INIT_17 = 256'h001A00722900000F001A00710D00003F001A00711200000F001A00717C00005F,
    pm.ram30_37.INIT_18 = 256'h001A00770800008F001A00731600006F001A00729100001F001A0072940000DF,
    pm.ram30_37.INIT_19 = 256'h001A00781200000F001A00787C00005F001A00780900000F001A00770C0000BF,
    pm.ram30_37.INIT_1A = 256'h001A00799100001F001A00799400006F001A00792900000F001A00780D00003F,
    pm.ram30_37.INIT_1B = 256'h001A00810800008F001A007D9500003F001A007C950000CF001A007A1600006F,
    pm.ram30_37.INIT_1C = 256'h001A00880800008F001A00819600007F001A00819600004F001A00810C0000BF,
    pm.ram30_37.INIT_1D = 256'h001A00981200000F001A00890E0000BF001A00890800008F001A00880E0000DF,
    pm.ram30_37.INIT_1E = 256'h001A00981200000F001A00981700004F001A00981200000F001A00981700000F,
    pm.ram30_37.INIT_1F = 256'h001A0099110000EF001A0099220000DF001A0099320000EF001A00986700009F,
    pm.ram30_37.INIT_20 = 256'h001A009F0C0000BF001A009F0800008F001A009F970000BF001A009B97000023,
    pm.ram30_37.INIT_21 = 256'h001A00B3970000BF001A00A1970000CA001A009F2300005F001A009F1600008F,
    pm.ram30_37.INIT_22 = 256'h001A00B49800001F001A00B49600009F001A00B4110000EF001A00B46E0000BF,
    pm.ram30_37.INIT_23 = 256'h001A00B70600007F001A00B70C0000BF001A00B7180000AF001A00B70600007F,
    pm.ram30_37.INIT_24 = 256'h001A00B70800002F001A00B70E0000DF001A00B7070000EF001A00B70D00005F,
    pm.ram30_37.INIT_25 = 256'h001A00BB0400004F001A00BB0C0000BF001A00BB0500003F001A00B70E0000DF,
    pm.ram30_37.INIT_26 = 256'h001A00BD9700009F001A00BD2000008F001A00BD9800005F001A00BC9800009F,
    pm.ram30_37.INIT_27 = 256'h001A00BE0400006F001A00BE0C0000BF001A00BE0500001F001A00BD2300005F,
    pm.ram30_37.INIT_28 = 256'h001A00CB0E00002F001A00CB0800000F001A00CA1500004F001A00BE9800003F,
    pm.ram30_37.INIT_29 = 256'h001A00CB0D00005F001A00CB0800002F001A00CB0D00005F001A00CB0A0000DF,
    pm.ram30_37.INIT_2A = 256'h001A00CB0D00005F001A00CB0800004F001A00CB0D00005F001A00CB070000EF,
    pm.ram30_37.INIT_2B = 256'h001A00CE0E00005F001A00CE0600005F001A00CB0E00002F001A00CB0600005F,
    pm.ram30_37.INIT_2C = 256'h001A00CE0C0000BF001A00CE070000EF001A00CE0C0000BF001A00CE0800004F,
    pm.ram30_37.INIT_2D = 256'h001A00CE0C0000BF001A00CE0A0000DF001A00CE0C0000BF001A00CE0800002F,
    pm.ram30_37.INIT_2E = 256'h001A00D70C0000BF001A00D70600007F001A00CE0E00005F001A00CE0800000F,
    pm.ram30_37.INIT_2F = 256'h001A00D72700000F001A00D71B0000FF001A00D70C0000BF001A00D70800004F,
    pm.ram30_37.INIT_30 = 256'h001A00D80C0000BF001A00D80600005F001A00D7260000AF001A00D7220000DF,
    pm.ram30_37.INIT_31 = 256'h001A00D86100002F001A00D8220000DF001A00D82A00007F001A00D81200002F,
    pm.ram30_37.INIT_32 = 256'h001A00DC0E00002F001A00DC0600005F001A00DB100000CF001A00DB9A00003F,
    pm.ram30_37.INIT_33 = 256'h001A00DC0E0000DF001A00DC0A0000DF001A00DC0E0000DF001A00DC0800004F,
    pm.ram30_37.INIT_34 = 256'h001A00DC0D00005F001A00DC070000EF001A00DC0E0000DF001A00DC0800002F,
    pm.ram30_37.INIT_35 = 256'h001A00DE2300005F001A00DE1200000F001A00DD2000008F001A00DD9600009F,
    pm.ram30_37.INIT_36 = 256'h001A00DF110000EF001A00DF9900006F001A00DF100000FF001A00DE9A00009F,
    pm.ram30_37.INIT_37 = 256'h001A00F31600008F001A00F36E0000BF001A00F36C00008F001A00DF200000EF,
    pm.ram30_37.INIT_38 = 256'h001A00F60C0000BF001A00F60800004F001A00F60C0000BF001A00F60800002F,
    pm.ram30_37.INIT_39 = 256'h001A00F70C0000BF001A00F70600005F001A00F61300004F001A00F6130000CF,
    pm.ram30_37.INIT_3A = 256'h001A00FB1200006F001A00FB6D00003F001A00F70D00005F001A00F70800004F,
    pm.ram30_37.INIT_3B = 256'h001A00FC1B0000DF001A00FC7B0000AF001A00FB110000CF001A00FB2B00001F,
    pm.ram30_37.INIT_3C = 256'h001A00FF110000EF001A00FE1600008F001A00FE6E0000BF001A00FC020000CF,
    pm.ram30_37.INIT_3D = 256'h011A00061200006F011A00066D00003F011A00029C00009F011A00019C00009F,
    pm.ram30_37.INIT_3E = 256'h011A0007220000DF011A00077B0000AF011A0006110000CF011A00062B00001F,
    pm.ram30_37.INIT_3F = 256'h011A00092300005F011A0009220000DF011A00096D00003F011A0007020000CF;
defparam
    pm.ram38_3F.INIT_00 = 256'h011A000D9D00004F011A000B110000EF011A000A1600008F011A000A6E0000BF,
    pm.ram38_3F.INIT_01 = 256'h011A002C0A00006F011A002B0F00007F011A000E9D0000BF011A000E2300005F,
    pm.ram38_3F.INIT_02 = 256'h011A002C1400000F011A002C3700004F011A002C390000FF011A002C0C0000BF,
    pm.ram38_3F.INIT_03 = 256'h011A002D3700008F011A002D390000FF011A002D0C0000BF011A002D0A00006F,
    pm.ram38_3F.INIT_04 = 256'h011A002D0D00005F011A002D1700000F011A002D0D00009F011A002D1200004F,
    pm.ram38_3F.INIT_05 = 256'h011A00340C0000BF011A0034180000AF011A0034180000AF011A00340A00006F,
    pm.ram38_3F.INIT_06 = 256'h011A0037370000AF011A00370F00007F011A00346000007F011A0034370000AF,
    pm.ram38_3F.INIT_07 = 256'h001B002E0C0000BF001B002E9F00002E011A00370D00005F011A00371200002F,
    pm.ram38_3F.INIT_08 = 256'h001B00301500006F001B00309F00004F001B00301200000F001B002E0C0000BF,
    pm.ram38_3F.INIT_09 = 256'h001B00310C0000BF001B00319F00002E001B0031180000EF001B00311700000F,
    pm.ram38_3F.INIT_0A = 256'h001B00379F0000B8001B00312C00002F001B00310C0000BF001B0031130000CF,
    pm.ram38_3F.INIT_0B = 256'h001B0037140000CF001B00371200000F001B00379F00004F001B00370D00009F,
    pm.ram38_3F.INIT_0C = 256'h001B00389F0000B8001B00389F00006F001B0038190000CF001B00381200000F,
    pm.ram38_3F.INIT_0D = 256'h001B003A110000EF001B00392B00008F001B00399F0000B8001B00382B00008F,
    pm.ram38_3F.INIT_0E = 256'h001B004D1100007F001B003A2B00005F001B003A2900000F001B003A9F0000B8,
    pm.ram38_3F.INIT_0F = 256'h001B004D0F0000BF001B004D2B0000EF001B004D0F0000BF001B004D1B0000FF,
    pm.ram38_3F.INIT_10 = 256'h001B004E0F00001F001B004E0C0000BF001B004E9F00002E001B004D2B00008F,
    pm.ram38_3F.INIT_11 = 256'h001B004E1200000F001B004E180000AF001B004E130000CF001B004E180000EF,
    pm.ram38_3F.INIT_12 = 256'h001B004F2900000F001B004F0F0000BF001B004E1300000F001B004E0C0000BF,
    pm.ram38_3F.INIT_13 = 256'h001B004F1600008F001B004F2E00003F001B004F1200004F001B004F120000AF,
    pm.ram38_3F.INIT_14 = 256'h001B00500D00003F001B00500F00007F001B00502C00002F001B00500C0000BF,
    pm.ram38_3F.INIT_15 = 256'h001B0051020000CF001B00501B0000DF001B00501C00001F001B00502A00007F,
    pm.ram38_3F.INIT_16 = 256'h001B00540C0000BF001B00549F00002E001B00511B0000DF001B00510F00007F,
    pm.ram38_3F.INIT_17 = 256'h001B0054130000CF001B0054180000EF001B00541700000F001B00540F00001F,
    pm.ram38_3F.INIT_18 = 256'h001B0056180000EF001B00560F00001F001B00560C0000BF001B00569F00002E,
    pm.ram38_3F.INIT_19 = 256'h001B00570C0000BF001B00571200000F001B0057180000AF001B0056130000CF,
    pm.ram38_3F.INIT_1A = 256'h001B0057220000DF001B00572C00002F001B00572300005F001B00571300000F,
    pm.ram38_3F.INIT_1B = 256'h001B00670C0000BF001B00670600009F001B0059A300000F001B0057110000EF,
    pm.ram38_3F.INIT_1C = 256'h001B0068140000EF001B00680D00003F001B00681200004F001B00670F00009F,
    pm.ram38_3F.INIT_1D = 256'h001B00691200004F001B00682A00007F001B00680F00009F001B00681200000F,
    pm.ram38_3F.INIT_1E = 256'h001B0069610000CF001B0069140000EF001B00691300006F001B00690C0000FF,
    pm.ram38_3F.INIT_1F = 256'h001B006A1B0000DF001B006A8A00006F001B006A1C00001F001B00692A00007F,
    pm.ram38_3F.INIT_20 = 256'h001B006B0F00007F001B006A1400002F001B006A0F00007F001B006A110000EF,
    pm.ram38_3F.INIT_21 = 256'h001B006E1200000F001B006E1200000F001B006B0D00005F001B006B0600009F,
    pm.ram38_3F.INIT_22 = 256'h001B006E0F00009F001B006E0D00003F001B006E1200004F001B006E110000EF,
    pm.ram38_3F.INIT_23 = 256'h001C00161B0000FF001C00160F00009F001B006E0F00007F001B006E2A00007F,
    pm.ram38_3F.INIT_24 = 256'h001C00171C00001F001C00171300000F001C00162B00001F001C00160F0000BF,
    pm.ram38_3F.INIT_25 = 256'h001C00181B0000DF001C00180F00007F001C00172A00007F001C00171B0000DF,
    pm.ram38_3F.INIT_26 = 256'h001C001B1400000F001C001B110000CF001C001BA5000059001C001B1B0000FF,
    pm.ram38_3F.INIT_27 = 256'h001C001E2C00002F001C001E1200000F001C001B150000AF001C001B1700002F,
    pm.ram38_3F.INIT_28 = 256'h001C001E1500004F001C001E1B0000FF001C001E1700002F001C001E130000CF,
    pm.ram38_3F.INIT_29 = 256'h001C001F140000EF001C001F0D00003F001C001F1700002F001C001F1200000F,
    pm.ram38_3F.INIT_2A = 256'h001C0023A5000059001C00201B0000DF001C001F0D00009F001C001F1200004F,
    pm.ram38_3F.INIT_2B = 256'h001C00392900000F001C0039A60000FF001C0039110000EF001C0023150000AF,
    pm.ram38_3F.INIT_2C = 256'h001C00391600008F001C00392E00003F001C00391200004F001C00391200002F,
    pm.ram38_3F.INIT_2D = 256'h001C003D1200000F001C003CA800001F001C003C2C00002F001C003C1200000F,
    pm.ram38_3F.INIT_2E = 256'h001C003D2A00007F001C003D0D00003F001C003DA60000FF001C003D2C00002F,
    pm.ram38_3F.INIT_2F = 256'h001C003E2D00001F001C003E2C0000BF001C003E1200006F001C003E1200006F,
    pm.ram38_3F.INIT_30 = 256'h001C0042140000EF001C00420D00003F001C00421200004F001C003F2C00002F,
    pm.ram38_3F.INIT_31 = 256'h001C00432B0000EF001C00430B00002F001C00432900000F001C0043A60000FF,
    pm.ram38_3F.INIT_32 = 256'h001C00450B00002F001C00442B00008F001C00440B00002F001C00442A00007F,
    pm.ram38_3F.INIT_33 = 256'h001C0051130000CF001C00511B0000FF001C00500F00009F001C00452900000F,
    pm.ram38_3F.INIT_34 = 256'h001C00511B0000DF001C0051140000EF001C00510D00003F001C00511700002F,
    pm.ram38_3F.INIT_35 = 256'h001C00521200004F001C0051020000CF001C00510D00009F001C00510F00007F,
    pm.ram38_3F.INIT_36 = 256'h001C00522C0000BF001C00520F00007F001C0052140000EF001C00520D00003F,
    pm.ram38_3F.INIT_37 = 256'h001C0053110000EF001C00534D00007F001C00530F0000BF001C0052020000CF,
    pm.ram38_3F.INIT_38 = 256'h001C00541200004F001C00541B0000FF001C00532D00001F001C00530F0000BF,
    pm.ram38_3F.INIT_39 = 256'h001C00552E00003F001C00551200004F001C00550F0000BF001C00540F00009F,
    pm.ram38_3F.INIT_3A = 256'h001C00561200004F001C00560F00007F001C00552A00007F001C00551600008F,
    pm.ram38_3F.INIT_3B = 256'h001C0056A600002A001C00560F0000BF001C00561600008F001C00562E00003F,
    pm.ram38_3F.INIT_3C = 256'h001C00571E00008F001C00571C00004F001C00571C00001F001C00562A00007F,
    pm.ram38_3F.INIT_3D = 256'h001C005CA60000BF001C005C1B0000FF001C00572D00001F001C00570F00007F,
    pm.ram38_3F.INIT_3E = 256'h001C005D0B00002F001C005C020000EF001C005C110000CF001C005C2B00001F,
    pm.ram38_3F.INIT_3F = 256'h001C005D0B00002F001C005D2900000F001C005DAB00007F001C005D2B0000EF;

endmodule
