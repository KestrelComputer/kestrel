`timescale 1ns / 1ps
module VRAM(
	input					RST_I,
	input					CLK_I,
	input		[12:0]	VF_ADR_I,
	input					VF_CYC_I,
	input					VF_STB_I,
	output				VF_ACK_O,
	output	[15:0]	VF_DAT_O,
	input		[12:0]	CPU_ADR_I,
	input		[15:0]	CPU_DAT_I,
	output	[15:0]	CPU_DAT_O,
	input					CPU_STB_I,
	output				CPU_ACK_O,
	input					CPU_WE_I
);

	reg				raw_ack;
	reg				ram_ack;
	wire	[15:0]	dat0, dat1, dat2, dat3, dat4, dat5, dat6, dat7;
	wire	[15:0]	cpu_dat0, cpu_dat1, cpu_dat2, cpu_dat3, cpu_dat4, cpu_dat5, cpu_dat6, cpu_dat7;
	reg	[15:0]	ram_q;
	reg	[15:0]	cpu_ram_q;
	reg				cpu_ram_ack;
	reg				cpu_raw_ack;

	assign	VF_ACK_O	= ram_ack;
	assign	VF_DAT_O = ram_q;
	assign	CPU_ACK_O = cpu_ram_ack;
	assign	CPU_DAT_O = cpu_ram_q;

	always @(*) begin
		ram_ack <= raw_ack & VF_CYC_I & VF_STB_I;
		cpu_ram_ack <= cpu_raw_ack & CPU_STB_I;

		case(VF_ADR_I[12:10])
			0:	ram_q <= dat0;
			1: ram_q <= dat1;
			2:	ram_q <= dat2;
			3:	ram_q <= dat3;
			4:	ram_q <= dat4;
			5: ram_q <= dat5;
			6:	ram_q <= dat6;
			7:	ram_q <= dat7;
		endcase

		case(CPU_ADR_I[12:10])
			0:	cpu_ram_q <= cpu_dat0;
			1: cpu_ram_q <= cpu_dat1;
			2:	cpu_ram_q <= cpu_dat2;
			3:	cpu_ram_q <= cpu_dat3;
			4:	cpu_ram_q <= cpu_dat4;
			5: cpu_ram_q <= cpu_dat5;
			6:	cpu_ram_q <= cpu_dat6;
			7:	cpu_ram_q <= cpu_dat7;
		endcase
	end

	always @(posedge CLK_I) begin
		raw_ack <= VF_STB_I & !raw_ack;
		cpu_raw_ack <= CPU_STB_I & !cpu_raw_ack;
	end

	wire vf_ram_0 = VF_ADR_I[12:10] == 0;
	wire vf_ram_1 = VF_ADR_I[12:10] == 1;
	wire vf_ram_2 = VF_ADR_I[12:10] == 2;
	wire vf_ram_3 = VF_ADR_I[12:10] == 3;
	wire vf_ram_4 = VF_ADR_I[12:10] == 4;
	wire vf_ram_5 = VF_ADR_I[12:10] == 5;
	wire vf_ram_6 = VF_ADR_I[12:10] == 6;
	wire vf_ram_7 = VF_ADR_I[12:10] == 7;

	wire cpu_ram_0 = CPU_ADR_I[12:10] == 0;
	wire cpu_ram_1 = CPU_ADR_I[12:10] == 1;
	wire cpu_ram_2 = CPU_ADR_I[12:10] == 2;
	wire cpu_ram_3 = CPU_ADR_I[12:10] == 3;
	wire cpu_ram_4 = CPU_ADR_I[12:10] == 4;
	wire cpu_ram_5 = CPU_ADR_I[12:10] == 5;
	wire cpu_ram_6 = CPU_ADR_I[12:10] == 6;
	wire cpu_ram_7 = CPU_ADR_I[12:10] == 7;

	RAMB16_S18_S18 r0(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_0),				.ENB(cpu_ram_0),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat0),						.DOB(cpu_dat0),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);

	RAMB16_S18_S18 r1(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_1),				.ENB(cpu_ram_1),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat1),						.DOB(cpu_dat1),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);

	RAMB16_S18_S18 r2(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_2),				.ENB(cpu_ram_2),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat2),						.DOB(cpu_dat2),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);

	RAMB16_S18_S18 r3(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_3),				.ENB(cpu_ram_3),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat3),						.DOB(cpu_dat3),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);

	RAMB16_S18_S18 r4(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_4),				.ENB(cpu_ram_4),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat4),						.DOB(cpu_dat4),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);

	RAMB16_S18_S18 r5(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_5),				.ENB(cpu_ram_5),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat5),						.DOB(cpu_dat5),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);

	RAMB16_S18_S18 r6(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_6),				.ENB(cpu_ram_6),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat6),						.DOB(cpu_dat6),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);

	RAMB16_S18_S18 r7(
		.WEA(1'b0),						.WEB(CPU_WE_I),
		.ENA(vf_ram_7),				.ENB(cpu_ram_7),
		.SSRA(RST_I),					.SSRB(RST_I),
		.CLKA(CLK_I),					.CLKB(CLK_I),
		.ADDRA(VF_ADR_I[9:0]),		.ADDRB(CPU_ADR_I[9:0]),
		.DOA(dat7),						.DOB(cpu_dat7),
		.DIA(16'hFFFF),				.DIB(CPU_DAT_I),
		.DIPA(2'b11),					.DIPB(2'b11)
	);


	defparam
r0.INIT_3F = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_3E = 256'h55555555555555555555555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_3D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_3C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_3B = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_3A = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_39 = 256'h55555555555555555555000000000000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_38 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_37 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA000C228AF1C2,
r0.INIT_36 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_35 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_34 = 256'h55555555555555555555010C228A8882AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_33 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_32 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA019822FA8882,
r0.INIT_31 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_30 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_2F = 256'h55555555555555555555C1D82A53F082AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_2E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_2D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA21F02A528882,
r0.INIT_2C = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_2B = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_2A = 256'h5555555555555555555521FC36228882AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_29 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_28 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAC1F8A223F1CF,
r0.INIT_27 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_26 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_25 = 256'h5555555555555555555501F000000000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_24 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_23 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAE1E0A0FB7228,
r0.INIT_22 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_21 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_20 = 256'h5555555555555555555501C0A0828A28AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_1F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_1E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA0180A0820A28,
r0.INIT_1D = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_1C = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_1B = 256'h555555555555555555558100BC8373EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_1A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_19 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA0000A282822A,
r0.INIT_18 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_17 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_16 = 256'h555555555555555555550000A282894DAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_15 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_14 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAE000BC837088,
r0.INIT_13 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_12 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_11 = 256'h55555555555555555555000000000000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_10 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_0F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAEF88088B8BE7,
r0.INIT_0E = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_0D = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_0C = 256'h55555555555555555555080088929208AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_0B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_0A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA080888A2A200,
r0.INIT_09 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_08 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_07 = 256'h55555555555555555555880808F3C387AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_06 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_05 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA081C088AA208,
r0.INIT_04 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_03 = 256'h5555555555555555555555555555555555555555555555555555555555555555,
r0.INIT_02 = 256'h55555555555555555555081C888A9208AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_01 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
r0.INIT_00 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAE8083EF38BE7;

endmodule
