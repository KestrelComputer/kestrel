`ifndef SIA_VH
`define SIA_VH

`define SIA_ADR_CONFIG		(0)
`define SIA_ADR_STATUS		(1)
`define SIA_ADR_INTENA		(2)
`define SIA_ADR_TRXDAT		(3)
`define SIA_ADR_zero0		(4)
`define SIA_ADR_zero1		(5)
`define SIA_ADR_BITRATL		(6)
`define SIA_ADR_BITRATH		(7)

`endif
