`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,

	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO,
	
	// SD Card Interface
	output			N2_SD_CLK_O,
	output			N2_SD_MOSI_O,
	output			N2_SD_CS_O,
	output			N2_SD_LED_O,

	input				N2_SD_MISO_I,
	input				N2_SD_WP_I,
	input				N2_SD_CD_I
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				gpia_ack_o;
	wire	[15:0]	gpia_dat_o;
	wire				gpia_stb_i;
	wire	[15:0]	gpia_port_o;

	assign N2_SD_CLK_O	= gpia_port_o[3];
	assign N2_SD_MOSI_O	= gpia_port_o[2];
	assign N2_SD_CS_O		= gpia_port_o[1];
	assign N2_SD_LED_O	= gpia_port_o[0];

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB00);		// B000-B003 : KIA
	assign gpia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB01);		// B010-B013 : GPIA 
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i & ~gpia_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	wire	[15:0]	gpia_mask			= {16{gpia_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)} | (gpia_mask & gpia_dat_o);
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | (gpia_stb_i & gpia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	GPIA gpia(
		.RST_I(N2_BTN0_I),
		.CLK_I(mgia_25mhz_o),
		.ADR_I(cpu_adr_o[1]),
		.CYC_I(cpu_cyc_o),
		.STB_I(gpia_stb_i),
		.WE_I(cpu_we_o),
		.DAT_I(cpu_dat_o),
		.DAT_O(gpia_dat_o),
		.ACK_O(gpia_ack_o),
		.PORT_I({13'h0000, N2_SD_MISO_I, N2_SD_WP_I, N2_SD_CD_I}),
		.PORT_O(gpia_port_o)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h03ABABAB03FF0000000000000000000000000000000000000000B800DA001E00,
progmem.ram00.INIT_01 = 256'h0D1015740000FF6BCB8BCB6BF303030303ABABAB03FFFF0B0B0B0B0BF3030303,
progmem.ram00.INIT_02 = 256'h15B8000000A41212F71215A4000094E00C101594000084E003101584000074E0,
progmem.ram00.INIT_03 = 256'hBA00E0F4000000E01212081216E0000000CC1212FD1215CC000000B81212FB12,
progmem.ram00.INIT_04 = 256'hFF141434000024E00410152400000E2E121261CE1AE00E000000F41212041216,
progmem.ram00.INIT_05 = 256'h000066E03678E014033066000050E03662E014E83050000034E03A4C1E141412,
progmem.ram00.INIT_06 = 256'hC2E0802415B0000092E0BAACE092E0F6A2E0A6009200007CE0E28EE06888E07C,
progmem.ram00.INIT_07 = 256'hB200E0B2FAE0B2F4E0B2EEE0B2E8E0DC000000B024B124241A7ECEE07EC8E094,
progmem.ram00.INIT_08 = 256'h000016E0DE38E0242E1BDE2CE02400012E4A160000DCE0B212E0B20CE0B206E0,
progmem.ram00.INIT_09 = 256'hFFB07600003CE0DE72E0241F1B1866E02E2013185AE02E2213DE4EE0241E1B3C,
progmem.ram00.INIT_0A = 256'h30003192161E16FF247EAEE07EA8E0BA00269EE0C416178C000076E0DE88E024,
progmem.ram00.INIT_0B = 256'hEAE0D0FCE03EF6E0EA0000CEE08EE6E0F6E0E0160030CE0000008C300131008C,
progmem.ram00.INIT_0C = 256'h12243EE032000022E0012615220000000E0112021AE00E000000003012000000,
progmem.ram00.INIT_0D = 256'h15780000006A26126A0000005601124862E056000046E0042615460000003201,
progmem.ram00.INIT_0E = 256'hBA000088E07EB6E07EB0E025011B25AA1A269EE025B025251A88000078E00028,
progmem.ram00.INIT_0F = 256'hBAE026251B8AF6E08AF0E08AEAE08AE4E08ADEE08AD8E08AD2E08ACCE02500B0,
progmem.ram00.INIT_10 = 256'h00E08A3CE08A36E08A30E08A2AE08A24E08A1EE08A18E08A12E02500B0000000,
progmem.ram00.INIT_11 = 256'h13427EE0282C134272E066000040E02C251B025CE000012C2511024CE0400000,
progmem.ram00.INIT_12 = 256'h0000ACE08AB8E0AC000088E068A8E00088A2127C2615BC94E088000066E02A2C,
progmem.ram00.INIT_13 = 256'h30F80000BCE000C23231FF3221180141181A31011A211A251202CEE0F43217BC,
progmem.ram00.INIT_14 = 256'h42E0103CE03000000EE01400000E2812FF2516021AE00E0000F8E0BE0AE03200,
progmem.ram00.INIT_15 = 256'h120020003170000052E0326CE0005266126C5EE052000030E0024EE00248E0FA,
progmem.ram00.INIT_16 = 256'h10C0E0BCBAE0BA0010B0E0ECAAE01F95B0729EE01E40B0CE92E0860000007022,
progmem.ram00.INIT_17 = 256'hE010FEE0BCF8E0F80010EEE0ECE8E072E2E01E41B0CED6E0CA000086E078C6E0,
progmem.ram00.INIT_18 = 256'h1040E0AE3AE03A001030E0EC2AE020007220E01E48B0CE14E0080000CAE07804,
progmem.ram00.INIT_19 = 256'hE0BC7EE07E001074E0EC6EE00022002011001E50B1CE56E04A000008E07846E0,
progmem.ram00.INIT_1A = 256'hC2E0C80010B8E0ECB2E0201C1372A6E01E51B0CE9AE08E00004AE0788AE01084,
progmem.ram00.INIT_1B = 256'h060010FCE0ECF6E072F0E01E77B0CEE4E0D800008EE078D4E010CEE054C8E0BC,
progmem.ram00.INIT_1C = 256'hE0DA3EE032000016002E0016002C119622E0160000D8E07812E0100CE0BC06E0,
progmem.ram00.INIT_1D = 256'h32E0787CE01076E0BC70E070001066E0EC60E000200022111850E01E69B0CE44,
progmem.ram00.INIT_1E = 256'h0080E078BAE010B4E08AAEE0AE0010A4E0EC9EE07298E01E7AB0CE8CE0800000,
progmem.ram00.INIT_1F = 256'h7E00E07EFAE07EF4E07EEEE07EE8E07EE2E07EDCE07ED6E07ED0E07ECAE0BE00,
progmem.ram00.INIT_20 = 256'h0004E0C03AE0C034E0C02EE0C028E0C022E0C01CE0C016E0C010E0040000BEE0,
progmem.ram00.INIT_21 = 256'h11001A003170000000600E01316000003EE0065CE01056E0F650E0A64AE03E00,
progmem.ram00.INIT_22 = 256'hE0CE0002BAE04CB4E09EE0AE0E179E000070E0909AE01C1213908EE0001C0018,
progmem.ram00.INIT_23 = 256'h31F8000000E8120031E800009EE00E013062DEE0E4006CD4E0009E0E013162C4,
progmem.ram00.INIT_24 = 256'h6240E04A000236E08230E02400000EE0EA20E01004300E000000F81212011008,
progmem.ram00.INIT_25 = 256'hE0107EE024E0FA74E078007A6AE000240E0131625AE064006C50E000240E0131,
progmem.ram00.INIT_26 = 256'hCA00011016B0000082E026ACE082E0EAA2E0A6008698E082E0920E1782000024,
progmem.ram00.INIT_27 = 256'h00D4E000D40E013162F0E0FA0002E6E0B2E0E0D40000B0E0CCD0E0B0E034C6E0,
progmem.ram00.INIT_28 = 256'h42E0003CE026E0360E172600000012A21201A21412000000FEA01201A014FE00,
progmem.ram00.INIT_29 = 256'h0EA131627AE084007670E000260EF1316A0C171096124854E0D64EE01448E052,
progmem.ram00.INIT_2A = 256'h000026E00E013062B2E0B8006CA8E02CA21E249CE02CE010019611868AE00026,
progmem.ram00.INIT_2B = 256'h013062FCE0020048F2E000BC0E013162E2E0EC0002D8E082D2E0BCE0CC0E17BC,
progmem.ram00.INIT_2C = 256'h00023EE00A38E022E0320E17220000060C2E0006031C114812E0060000BCE00E,
progmem.ram00.INIT_2D = 256'h0131627CE086000272E0886CE0600000002210120858E000220E01316248E052,
progmem.ram00.INIT_2E = 256'h0026BEE040B8E00E0000100031A0000060E00E01306296E09C00348CE000600E,
progmem.ram00.INIT_2F = 256'hFA000000A00EFF3162F0E0A0E0A0E6E084E0E028DAE0BED4E024CEE062C8E0EA,
progmem.ram00.INIT_30 = 256'h1A121C1A213000001CE0FC2CE01C001C0000FAE0001C1E021C141C0023181C17,
progmem.ram00.INIT_31 = 256'h82E076000054E03272E0326CE03266E03260E054000000301C12501C141A0213,
progmem.ram00.INIT_32 = 256'hAE0112011015AE000098E078AAE01C363098000076E05694E0568EE05688E056,
progmem.ram00.INIT_33 = 256'h0600B0FCE0F0000000D61212011216C4E2E0D6000000C21212FE1215C2000000,
progmem.ram00.INIT_34 = 256'h42E0C43CE03000000EE0F22CE09A26E01A3430C41AE00E0000F0E0F6000406E0,
progmem.ram00.INIT_35 = 256'h1080E0327AE00874E00EAA30740017187A12B05CE07256E04A000030E000001E,
progmem.ram00.INIT_36 = 256'hC2E0B6000084E010B2E08A0052FF1B26021A26001A0EAC12B090E08400004AE0,
progmem.ram00.INIT_37 = 256'h0C110E1212B0F6E0A2F0E01EEAE0D8E4E0D80000B6E086D4E09ACEE01A5430C4,
progmem.ram00.INIT_38 = 256'hE0103EE00438E03800B02EE01E28E01C0000D8E01018E04C12E0080CE0000ECC,
progmem.ram00.INIT_39 = 256'h000000000000000000000000000000000000000000000000000000000000001C,
progmem.ram00.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'hC8CA6232180F00000000000095000000000000000000000000000D1E0D1E0E1E,
progmem.ram01.INIT_01 = 256'h000012001300FFD6D3D1D3D6CFC0C0C8C8CA6232180FFFD0D0D0D0D0CFC0C0C8,
progmem.ram01.INIT_02 = 256'h12001300E000B013FFB012001300001200001200130000120000120013000012,
progmem.ram01.INIT_03 = 256'h000111001300E000B01300B012001300E000B013FFB012001300E000B013FFB0,
progmem.ram01.INIT_04 = 256'hFF0012011300011200B0120113000131B0B012000111011300E000B01300B012,
progmem.ram01.INIT_05 = 256'h1300011201011100001101130001120101110003110113000112010117000013,
progmem.ram01.INIT_06 = 256'h011100001A011300011200011101120001110117011300011200011101011101,
progmem.ram01.INIT_07 = 256'h0102110101110101110101110101110113002E01004100001A01011101011101,
progmem.ram01.INIT_08 = 256'h1300021201021100001A010211001B0000110213000112010211010211010211,
progmem.ram01.INIT_09 = 256'h0011021300021201021100001A02021100001202021100001201021100001A02,
progmem.ram01.INIT_0A = 256'h00001102001300FF110102110102110217010211020012021300021201021100,
progmem.ram01.INIT_0B = 256'h021202021102021102130002120202110002110020110213002E020000112E02,
progmem.ram01.INIT_0C = 256'h16030311031300031200001A031300E0030016030311031300E0030012031300,
progmem.ram01.INIT_0D = 256'h12031300E003001A031300E0030016030311031300031200001A031300E00300,
progmem.ram01.INIT_0E = 256'h0313000312010311010311000016000317010311004100001A03130003124000,
progmem.ram01.INIT_0F = 256'h031200001A030311030311030311030311030311030311030311030311000011,
progmem.ram01.INIT_10 = 256'h0412030411030411030411030411030411030411030411030411000011041300,
progmem.ram01.INIT_11 = 256'h12040411000012040411041300041200001A0404114B0000001A040411041300,
progmem.ram01.INIT_12 = 256'h130004120404110413000412040411E004041700001A03041104130004120000,
progmem.ram01.INIT_13 = 256'h110413000412E0040041FF00310000210000410000B100001A04041104001204,
progmem.ram01.INIT_14 = 256'h05110505110513000512051EE005051700001A04051105130004120405110002,
progmem.ram01.INIT_15 = 256'h13000000110513000512050511E0050517030511051300051204051104051104,
progmem.ram01.INIT_16 = 256'h0105110305110517030511020511000011050511000011000511051300E00500,
progmem.ram01.INIT_17 = 256'h1101051103051105170305110205110505110000110005110513000512020511,
progmem.ram01.INIT_18 = 256'h0106110406110617030611020611001305061100001100061106130005120206,
progmem.ram01.INIT_19 = 256'h1103061106170306110206113000000013020000110006110613000612020611,
progmem.ram01.INIT_1A = 256'h0611061703061102061100001205061100001100061106130006120206110106,
progmem.ram01.INIT_1B = 256'h0717030611020611050611000011000611061300061202061101061105061103,
progmem.ram01.INIT_1C = 256'h110607110713000700112E074007170007110713000612020711010711030711,
progmem.ram01.INIT_1D = 256'h0712020711010711030711071703071102071130000000130707110000110007,
progmem.ram01.INIT_1E = 256'h0007120207110107110407110717030711020711050711000011000711071300,
progmem.ram01.INIT_1F = 256'h0108110107110107110107110107110107110107110107110107110107110713,
progmem.ram01.INIT_20 = 256'h0008120708110708110708110708110708110708110708110708110813000712,
progmem.ram01.INIT_21 = 256'h130000C0110813002E0800001108130008120808110108110008110008110813,
progmem.ram01.INIT_22 = 256'h1108170308110608110812080012081300081206081100001206081130000000,
progmem.ram01.INIT_23 = 256'h110813002E08000211081300081200A01108081108170308112E080080110808,
progmem.ram01.INIT_24 = 256'h08091109170309110709110913000912080911000011091300E0080013000000,
progmem.ram01.INIT_25 = 256'h12090911091208091109170309112E0900E01108091109170309112E09008011,
progmem.ram01.INIT_26 = 256'h0917000012091300091209091109120809110917000911091209001209130009,
progmem.ram01.INIT_27 = 256'h0009122E09008011080911091703091109091109130009120509110912070911,
progmem.ram01.INIT_28 = 256'h0A110A0A110A120A00120A1300E00AC01300C0120A1300E009C01300C0120913,
progmem.ram01.INIT_29 = 256'h009811080A110A17000A112E0A0098110A0015000A17030A11090A110A0A1101,
progmem.ram01.INIT_2A = 256'h13000A12009811080A110A17030A110A0A17030A110A3100000A17000A112E0A,
progmem.ram01.INIT_2B = 256'h0C11080A110B17030A112E0A008011080A110A17030A11070A110A120A00120A,
progmem.ram01.INIT_2C = 256'h17030B11060B110B120B00120B13000B00112E0B000B17030B110B13000A1200,
progmem.ram01.INIT_2D = 256'h8011080B110B17030B11050B110B1300E00B00130B0B112E0B008011080B110B,
progmem.ram01.INIT_2E = 256'h17010B11080B110013000000110B13000B1200FF11080B110B17030B112E0B00,
progmem.ram01.INIT_2F = 256'h0B13002E0B000011080B110B12080B11090B110A0B110A0B110B0B110B0B110B,
progmem.ram01.INIT_30 = 256'h00230000120C13000C120B0C1100130C13000B120C00130000120000110C0012,
progmem.ram01.INIT_31 = 256'h0C110C13000C120C0C110C0C110C0C110C0C110C1300E00C0013000012000014,
progmem.ram01.INIT_32 = 256'h0C001600B0120C13000C120C0C1100D3110C13000C120C0C110C0C110C0C110C,
progmem.ram01.INIT_33 = 256'h0D170C0C110C1300E00CB01300B0120C0C110C1300E00CB013FFB0120C1300E0,
progmem.ram01.INIT_34 = 256'h0D110C0D110D13000D120C0D110C0D110000110C0D110D13000C120C1E000D11,
progmem.ram01.INIT_35 = 256'h0D0D110D0D11000D1100AA110D0416000D170C0D11080D110D13000D12C01E0C,
progmem.ram01.INIT_36 = 256'h0D110D13000D120D0D110D1EC0FF1600C01B00C013000D170C0D110D13000D12,
progmem.ram01.INIT_37 = 256'h0E17000E170C0D110B0D110C0D110C0D110D13000D120D0D110C0D110000110C,
progmem.ram01.INIT_38 = 256'h120D0E11000E110E170C0E110C0E110E13000D120D0E110D0E11000E113000CC,
progmem.ram01.INIT_39 = 256'h000000000000000000000000000000000000000000000000000000000000000E,
progmem.ram01.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
