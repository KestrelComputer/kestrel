`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,
	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:12] == 4'b1011);	// B000-B001 : KIA (B002-BFFF = repeats)
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)};
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h41014671000141FF0A16010C1420000010E00A0C13100000000000000F00F400,
progmem.ram00.INIT_01 = 256'hFF0A1474000000640C00316400004AE00C000CFF24600C174A000020E0000C0C,
progmem.ram00.INIT_02 = 256'h00ACC0126C0E16AC000088E012A8E076A2E000889C12690E1688000000740C12,
progmem.ram00.INIT_03 = 256'h7D0E16F40000D0E012F0E022EAE000D0E4127A0E16D00000ACE012CCE066C6E0,
progmem.ram00.INIT_04 = 256'h0000002802120E021328000018E00A0613180000F4E01214E04C0EE000F40812,
progmem.ram00.INIT_05 = 256'hE08800F002166E000058E05E6A1E0100155800003CE002521B0E0E120002163C,
progmem.ram00.INIT_06 = 256'h021E9CE070B8E0BC00E002165AA8E09C00006EE03E98E05A92E002006EE02A84,
progmem.ram00.INIT_07 = 256'hE01AFEE0F20000C6E0CC008AEAE0AEE4E0D2DEE0F6D8E09ED2E0C600009CE0A2,
progmem.ram00.INIT_08 = 256'hFFBFBB17F2DC2F5FC5FE5FCB7EBFBF5F2FFFFFF89700F2E0C810E0120AE06604,
progmem.ram00.INIT_09 = 256'hFFFB9DFFBF7CFF5F9717B21797E52BFFFBFF2FFE5980FF22242FBFE55FF2FC5E,
progmem.ram00.INIT_0A = 256'hF1FDFFFEF7BE92229292922224FF7E7FDEFFD8FFEFB1FCFF97FEBFFF6596FEFB,
progmem.ram00.INIT_0B = 256'hFFFFFF162FFFF81DFFFDC2F8FB5E5DBEF9F7FBF1BBBFE2FFFFFFBEFFFFBFE2FF,
progmem.ram00.INIT_0C = 256'h972AFFFFFFFF6CFE2D2B7EFFFFC22CB216B2BFF8C003030E3BBFDFFCE000BF6E,
progmem.ram00.INIT_0D = 256'hFFCBC5C7FFFFFF5C92FFF2BFFFBFEF7EF0F87FBBBFBB5FC5BCE1FEFF241278FF,
progmem.ram00.INIT_0E = 256'h5F2D00000000200000000020BBFDC5FFE5E2EDE27EDF5FF95FC5FDFFFFFF7E2B,
progmem.ram00.INIT_0F = 256'hC57F8B26C4FEFFFBFFFFFFAF7FFFFFDDDFF1F7BDDF7FF2C5FFBFFB5FFD2FFF77,
progmem.ram00.INIT_10 = 256'hF88BF8FFFF24F0F9FFE73FF297FF3F4949F1F1912CBDFDF997FFBFDFC5F7FFFF,
progmem.ram00.INIT_11 = 256'hF9BFFFABCBFFBF8500000000000048F2FFBFFFE2592E9716E2FE7FE597F97E79,
progmem.ram00.INIT_12 = 256'hCC8CE5FCFFB6E2CB49FFD7D7FFF9FFFFFFFFF87F97F9FFFEFCFE5FE5FEFF7F5F,
progmem.ram00.INIT_13 = 256'h7BDFF97F5FFE2FFFEF6FF9FDF75BDF99F397D7E557FFFEFD5957E2FF97E6F1CC,
progmem.ram00.INIT_14 = 256'h5FFFF998F9FF77F77FFBFF2FFCDFF1F2FD7B7F25F8E5975F7CBFFFFFBF972FDB,
progmem.ram00.INIT_15 = 256'h5F92BEFF8BBEFFC55FF2CBFFFFC57FFDFCFF452FFCE225FCE2F9321244915FFF,
progmem.ram00.INIT_16 = 256'h49F75E0B4849249292CBF97FFD856619FDBF97FFFF655FCBBFDFFF17FFFFF97F,
progmem.ram00.INIT_17 = 256'hBFAF7C450402082021410410422110211020418108088484F8F876127D5B16CB,
progmem.ram00.INIT_18 = 256'h482FF2E7F2FFFFFBBFFFFFFFFFDFFFE5FFFEFF92ED7F725BFFAFF797FFF2FFFF,
progmem.ram00.INIT_19 = 256'hFFFFFF8BFBEFFFF917EDFAFBFFFEED7FFF7D95F8FFFF7F7F5F5FFFDE7FBB1624,
progmem.ram00.INIT_1A = 256'hFB7FEFFFF7FFF67FBFFFE5FB7EF22BE589FFFFAFFF77927FFBFBFFF7FFEF7D7D,
progmem.ram00.INIT_1B = 256'h0000209249248244BFFFF7FEDFFE7FAFFFFDFFFFFECBFF5FFFBFFEDF5BBFFFFF,
progmem.ram00.INIT_1C = 256'hE6FFFF5FF3FEFF3FE57FCFF95FF857FFFFC27F857EDFFFFBFFAF5FFF7FC27E08,
progmem.ram00.INIT_1D = 256'hFFDFFCF22FF8FFDBFFFFF1FFBFED8BFB5FE52FF2FEFF7FBCFFF7CBBE81F81244,
progmem.ram00.INIT_1E = 256'h85FFFFB51FFFFFF1FF62FFF1C28B8AFE7FFE7F6E25F7F7F2EFFFFFEFFFFFF7EF,
progmem.ram00.INIT_1F = 256'hDF77BB97FDC5EF7BF5B7FDDF7FAF7BEFEDEBFBF7F7DDEDF85FBFFFFFFF5FFC2F,
progmem.ram00.INIT_20 = 256'h9249247C97F9BFCBEC7B2FF8BFE2FBFFFF7717EE7FFFFFF8F71749775FB9F75F,
progmem.ram00.INIT_21 = 256'h0000000000000000000000000000000000000000005E2FFFAECA57DFFD544524,
progmem.ram00.INIT_22 = 256'hF7E5BFDFBBDBCB7BDDBBBFBFFB44F8FFF9FF2FF2F92400000000000000000000,
progmem.ram00.INIT_23 = 256'hFEB777EE2DFFFFFFFFFFFF5FFF2F7DDDDFEFF7FFFFE5FCFFBEBF2FEEEFDBDF65,
progmem.ram00.INIT_24 = 256'hFFEFFFFFE2FEFEFFFBF8FFF5BFFFFFFF8BFEFFFF498BFFE26F8924792E7BEDFB,
progmem.ram00.INIT_25 = 256'hBFE5CBFFFF97EFFF2FFFFFFFBF77EFF7EEFFC9E2577DFFDEFFC5F1FFFF7FFFF7,
progmem.ram00.INIT_26 = 256'hF7FCFFEFEFEFBEFB8BF7FFFFEFF897FFFFFFFFEFFFF6DFFFF6FBCAF7FF7FFF57,
progmem.ram00.INIT_27 = 256'h5FBCCAAF2FCBDFF8BF2CBEBF2F0BFFDFFFF6FFEFBAC5FF00000400107FEEFFFF,
progmem.ram00.INIT_28 = 256'hFFFE5B7F2FDF7E5F17EFFE78F9EFBB2BB9F7FFFFFFC5FFFF491222912489F9EE,
progmem.ram00.INIT_29 = 256'hFCDD17DFBF0A16E0807F24EF2BFCFCFFFFFEF2FDEFF67FBFBE77FDEE775EBFDD,
progmem.ram00.INIT_2A = 256'h492492492492492448F217C5FE77DFFFFE3BF7DFBFFFFDC5F77FDFBFDF775DFB,
progmem.ram00.INIT_2B = 256'h4992644924669992269249FFF75FFFFF22E8FDAFF2FF2F242492492466666692,
progmem.ram00.INIT_2C = 256'h4999922664249264996699264992494999922664242664494924266449492426,
progmem.ram00.INIT_2D = 256'hFF1FEFFFE5AFFEDFD7EF88F8AF32DC7FDF644999922664249292266449999249,
progmem.ram00.INIT_2E = 256'hDF7FADFDDFFFFF17FFFFCAFFFFF9FFFFDEFFFFFC24AFFFE5FF494491FE2EDFFF,
progmem.ram00.INIT_2F = 256'hCBF2F1D9FEFB5F78FF7FFBFFC6F67FFFFF090000000000000020894989922497,
progmem.ram00.INIT_30 = 256'h0000000000000000EFFFF1EFF7BEDFF7FDF7BECB3BFD7777777DFFE5EE972292,
progmem.ram00.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'h12000051800014FF00120000120013000012C00012001300000000000000011E,
progmem.ram01.INIT_01 = 256'hFF00120013002E000000110013000012001300FF110000120013000012300000,
progmem.ram01.INIT_02 = 256'hE00000170000120013000012000011000011E0000017000012001300E0000013,
progmem.ram01.INIT_03 = 256'h0000120013000012000011000011E00000170000120013000012000011000011,
progmem.ram01.INIT_04 = 256'h1300E001B01B00B01A01130001120000120113000012000111000111E0000117,
progmem.ram01.INIT_05 = 256'h11011700B01A011300011201011700B01A0113000112B0C01300001380B01A01,
progmem.ram01.INIT_06 = 256'hB01B0112010111011700B01A0101110113000112010111010111B01B01120101,
progmem.ram01.INIT_07 = 256'h110101110113000112011E000111000111000111000111010111011300011201,
progmem.ram01.INIT_08 = 256'hFEE5BC78EFBFFFE3FE1FC5FE5FE5FCBCDEFFFFBFE50001120102110002110002,
progmem.ram01.INIT_09 = 256'hCBBFFFFFE292F9F2E5FFC9FC2EFF9797FFEFF7577FFCF71724FCF7F897FCBF2F,
progmem.ram01.INIT_0A = 256'h7EF7FFF6AD2F484449442444916F2FFBF1E5BFFFBF6558FFFF5FFFFCFFDCDFF7,
progmem.ram01.INIT_0B = 256'hE1FF052FDF7FAFE58BFFFFBFFDFFF1FC7F17FF7DFEFDFCFBFFFFFFEDEFFEF517,
progmem.ram01.INIT_0C = 256'hFFEFFEFFFFFF2FF9FF9757EF2FC5B2CB2CCB2C031DBFBFFCF0C083010E772FF8,
progmem.ram01.INIT_0D = 256'h92FFEF7FFFDF975F49E4FFFF7FC5F300073B9DF7FFF38BFC5F63577F5E498959,
progmem.ram01.INIT_0E = 256'hFFDE01000000000100000000FFF7BE2FFFFFFFDF2FF9FB7ECB7CEFFDF8E25F7F,
progmem.ram01.INIT_0F = 256'hEFFFE12F0C2FBF7FBFFF8BFFF8F1C5F7BF7F7DC58B77EF7FDFFFF777FCBBFFE2,
progmem.ram01.INIT_10 = 256'h59FFBFFFF2BF7E7FE1E22FFEF39F2F7F24227B7D48FAF87FE5FFCBDCFBFF0BFF,
progmem.ram01.INIT_11 = 256'h7EFFFCFFFFFFF8FC25000000000082FC2ECBC5CB7FFCF35FFF5FE579957F5DF9,
progmem.ram01.INIT_12 = 256'hCCCCF9AF155FF8FF652EEBE5AF77FFF22FF2B297F97F97FF5D5FE5FE5FE5F2F9,
progmem.ram01.INIT_13 = 256'hBFBF77EFF7FEFEFFEFFE25FF7DBE127F2FFFCB752B2E5FFF2596FE97FF2F7FCB,
progmem.ram01.INIT_14 = 256'h95FCCBBF7FFFF7FCFFBFEFC5BFF27DEFFFCBFFF9B1F2CB2FBE99FCF7FD8A97F7,
progmem.ram01.INIT_15 = 256'hE1E9A578FFC4FFBFDFFEFFFFFFF7E7F1BF7BFEF2BEFB8B91F27FFF238922C8FC,
progmem.ram01.INIT_16 = 256'h6E24E2DC9324924944E07EC1D98B2E8C7FCB7FDFF7FFE6DEF7FFE2BFBDFF7BFF,
progmem.ram01.INIT_17 = 256'hFFCC24FF220812820804108210088408428208088044212088BF5F1689B1EC3B,
progmem.ram01.INIT_18 = 256'h919249C5FFFFFFDFFFFED6FF2FFFFAFFD717EF57FDFFB9E5FEC5FCE5FF4BD7DF,
progmem.ram01.INIT_19 = 256'hF1FFFFEFFFFF176FFFFFEFFFFF2FFFFAF9EFFFBFDEFBEDF9F1FCF9FFFBE52C89,
progmem.ram01.INIT_1A = 256'h7FDFCBDDF2DFFFCBF7FFFEFD5FFF77FF17FFFF729CE249BFF997FF7FBECAFFF1,
progmem.ram01.INIT_1B = 256'h000000492492242495C2FFFFDF2EFFFFF8FF7FDF2BCBFFDFFECB2496F29217BF,
progmem.ram01.INIT_1C = 256'h623FE5F3FE5F3FE5FFCFF97FF3B8C5BCE2BBFF7FFF85018B0BF7F8FCC5BF2FB1,
progmem.ram01.INIT_1D = 256'hBDEFB7FEFFAFFFFFC58B7FFFFFE2BEFDEBFCFFEC5D7ADEBFEFFF2FA2F8572F89,
progmem.ram01.INIT_1E = 256'hFE17FFBFF8FE9F5FFFF7FF7FFFFFFF5F9549CBF9B9997FE5FDFFEFFFFFEFFFFF,
progmem.ram01.INIT_1F = 256'hFDDFEFE5FFFBBF16F5FF5EBFFFD5D55DBAEFDFDEEBAFEFBFFFBCFCFFFFFFBC0B,
progmem.ram01.INIT_20 = 256'h492492BFF97FCBFCBFFF99BFFFFC17FF8BFFF1FFEEC5BBBF7FFF33F2EF71F8FB,
progmem.ram01.INIT_21 = 256'h0000000000000000000000000000000000000000004077EFF2FCDDF6EF975592,
progmem.ram01.INIT_22 = 256'hF9F2FFFDEFFDFFBFFB7FF7FC5F9722977FFFFF497DBF01000000000000000000,
progmem.ram01.INIT_23 = 256'h2E7FFBFFDFFEFFFFFFFF85FFF9FFBCF7777DDD62FBF25F17FBDBFDFFEDFEBDFF,
progmem.ram01.INIT_24 = 256'hCBF7FF9725FF2FFF2FBFFFFFDFD8FF8BF25FFFE222161DCEBF11887F5BBFF9BC,
progmem.ram01.INIT_25 = 256'hF6FFFFFFFFFFFDFFFFFFE5CB8BB8BF7EFBDF17DF7FFCFF2BFFFF57FFFFFFF1FF,
progmem.ram01.INIT_26 = 256'hFF5FFFFFFBBFFBEFBEFDFFFFFFBEFFFFFF62FF2FE22F65E257BFFF7E2FFFD9FF,
progmem.ram01.INIT_27 = 256'hF8BCF22BFC89BF5F7758EEBBF8FCFBFF0B17FFDDFFDE2F1200400000BFF1EEFF,
progmem.ram01.INIT_28 = 256'h5FDFBFFEC5BF2FBFBCDFB7BB7F778BF37EEFFBFEFF8BEFFF8A24491148127FF1,
progmem.ram01.INIT_29 = 256'h0FF77FEFDFBF0B7EF9C749F7BEBEBFCBCB77EF8BF6B5F7EBFBD7DEFB9649F6FF,
progmem.ram01.INIT_2A = 256'h249249249249249291FCCBFF2FFFBBFFCAFFFFBFFFE08BFFF8FD17C578FFF1F8,
progmem.ram01.INIT_2B = 256'h9966992692492664494924C6FFFFECFF22B1FFFEFCFFFE4C9249249249666666,
progmem.ram01.INIT_2C = 256'h9226644999924999264992649966249226644999924999922692499992269249,
progmem.ram01.INIT_2D = 256'hFFFFFFEFFF7EF7FFD7D725BFFFC55FE22F859226644999924964499992266424,
progmem.ram01.INIT_2E = 256'hDFDDFFFFEB7777CBCBFFF7FFFF7FFF2FFFFFFFBFB292FC7FFF2592225CFDFFEF,
progmem.ram01.INIT_2F = 256'hF7F7FB7FDFFEFEFCDF7FD97D5F2F7EDF176200000000000000001224244448DE,
progmem.ram01.INIT_30 = 256'h00000000000000007EBD6F75FE5FFBFFFFCB5FFBFFEFBBF7FFFFFFE55EE54449,
progmem.ram01.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
