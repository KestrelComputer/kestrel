`ifndef SIA_VH
`define SIA_VH

`define SIA_ADR_CONFIG		(0)
`define SIA_ADR_STATUS		(1)

`endif
