`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,
	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:12] == 4'b1011);	// B000-B001 : KIA (B002-BFFF = repeats)
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)};
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h000C3818660000000000000000000000000000000F0000000000000000000A00,
progmem.ram00.INIT_01 = 256'h00601C06603018007E66C67E7C7C666006667E787C3C2004003C1C0C3C180000,
progmem.ram00.INIT_02 = 256'h3828100010000000FF8080E0FFFF000000FF0208208036180000000800000018,
progmem.ram00.INIT_03 = 256'h1020002810102028083C28102070102010202E281020C03038007C0838103800,
progmem.ram00.INIT_04 = 256'h24186C3E660000000000000000000000000000000F0040280802281020481020,
progmem.ram00.INIT_05 = 256'h18603006601818600666C618666676600666606C6666300C1866301C66240000,
progmem.ram00.INIT_06 = 256'h1C001044380000007FC040E0FFFF00000000020820806C180000001800000018,
progmem.ram00.INIT_07 = 256'h2810000028082000104C00281048281028105800281020104400F41004287400,
progmem.ram00.INIT_08 = 256'h18306858240000000000000000000000000000000F004000103C002810302810,
progmem.ram00.INIT_09 = 256'h007C303E7C0C3C300C3C6C186666766006666066666E18181866603C06660000,
progmem.ram00.INIT_0A = 256'h64001038540007E03FE020E0FF000000FF000208208000187E66663C5E7C5C18,
progmem.ram00.INIT_0B = 256'h38386C383838380000543838384438387C7C58000000C4104400F40018106C7C,
progmem.ram00.INIT_0C = 256'h7E30323C000000000000000000000000000000000F005844444C383838080000,
progmem.ram00.INIT_0D = 256'h18667C6666003C1818186C187C7C7E60067E78667C6A0C30003C7C6C0C660000,
progmem.ram00.INIT_0E = 256'h3C000028500018181FF010E0FF00000000000208208000180C3C661860666618,
progmem.ram00.INIT_0F = 256'h44441204040424444454444444E4101040408C101010287C3800740020007404,
progmem.ram00.INIT_10 = 256'h18306C1A0000000000000000000000000000000F000064444454444444383030,
progmem.ram00.INIT_11 = 256'h186630666600660C303C381878606E6066666066666618180066667E30660010,
progmem.ram00.INIT_12 = 256'h7C001038540010080FF808E0000000FF000002082080001818183C1860666618,
progmem.ram00.INIT_13 = 256'h7C7C7E3C3C3C384444544444444410106070F8282828D408000014003C006C00,
progmem.ram00.INIT_14 = 256'h24186C7C0000000000000000000000000000000F000064444464444444441010,
progmem.ram00.INIT_15 = 256'h1866306666000006606638186C606E606666606C6660300C1866660C60241818,
progmem.ram00.INIT_16 = 256'h000010443800200407FC04E0000000000000020820800018303C3C18607C6618,
progmem.ram00.INIT_17 = 256'h404090444444204444644444444810104040884444442C287C00140000006C00,
progmem.ram00.INIT_18 = 256'h000C3A180000000000000000000000000000000F000058444478444444441010,
progmem.ram00.INIT_19 = 256'h1866303E7C0000007E6610186660667E3C6660787C3C2004183C3C0C7E181810,
progmem.ram00.INIT_1A = 256'h000010001000200403FE02E00000FF0000000208208000187E66180C6060660C,
progmem.ram00.INIT_1B = 256'h38386E3C3C3C203838783838387038387C7C8E7C7C7C5C380008140000003800,
progmem.ram00.INIT_1C = 256'h000000000000000000000000000000000000000F000040383880383838383838,
progmem.ram00.INIT_1D = 256'h7000000000000000000000000000000000000000000000000000000000000020,
progmem.ram00.INIT_1E = 256'h000000000000200401FF01E00000000000000208208000000000000000600000,
progmem.ram00.INIT_1F = 256'h0000000000000000000000000000000000000044444404080010000000000000,
progmem.ram00.INIT_20 = 256'h8000800080008000800080008000800080008000800040000000000000000000,
progmem.ram00.INIT_21 = 256'h0202020202010101010101010100000000000000004543413836343230008000,
progmem.ram00.INIT_22 = 256'h0606060606050505050505050504040404040404040303030303030303020202,
progmem.ram00.INIT_23 = 256'h0A0A0A0A0A090909090909090908080808080808080707070707070707060606,
progmem.ram00.INIT_24 = 256'h0E0E0E0E0E0D0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0A0A0A,
progmem.ram00.INIT_25 = 256'h0017800A1470000000560A12020A140A00235600000F0F0F0F0F0F0F0F0E0E0E,
progmem.ram00.INIT_26 = 256'hE01442121212AE000000900A12500A140A2BFF0AA190000070E076005888E08C,
progmem.ram00.INIT_27 = 256'h0000E2E0001200F811001215E2000000C2121831C2E0D80017E71214C20000AE,
progmem.ram00.INIT_28 = 256'h110010153200000012104F3112E0280017B01014120000FCE0C40EE0E408E0FC,
progmem.ram00.INIT_29 = 256'hB080E0011016FE74E04E6EE06200004CE0145EE03458E04C000032E000100048,
progmem.ram00.INIT_2A = 256'h9E0A12500A140C00130C120A0CA19E0000008A0C120814A48A0000622E0A0041,
progmem.ram00.INIT_2B = 256'h00C4FEE0020017800C14E6000000C20A12020A140C02130C120A0C21C2000000,
progmem.ram00.INIT_2C = 256'h3A000024E07236E00A003024000006E0E820E00C8013000A0031060000E6E0EC,
progmem.ram00.INIT_2D = 256'h7A00003AE09276E09270E0926AE09264E0925EE09258E09252E0924CE06446E0,
progmem.ram00.INIT_2E = 256'hA0C0E0A0BAE0A0B4E0A0AEE0A0A8E08CA2E0649CE0900000007A121200100031,
progmem.ram00.INIT_2F = 256'h13120812181216EC0000D6E072E8E008E2E0D6000090E0A0D2E0A0CCE0A0C6E0,
progmem.ram00.INIT_30 = 256'h104A124F10169234E02800000012100031EE1EE0120000ECE0D80EE0ECE01201,
progmem.ram00.INIT_31 = 256'h2A80E00820B06E000054E02A6AE008B046081454000028E01450E028E0100113,
progmem.ram00.INIT_32 = 256'h1BB800009EE056B4E008B05609149E000084E0569AE008000F09158400006EE0,
progmem.ram00.INIT_33 = 256'h00EC0612FF0614EC000000D80112010015D8000000B8021286D0E0A0CAE00902,
progmem.ram00.INIT_34 = 256'h00002E0E01312E000010012E10002E280617EE1CE01000000000060031000000,
progmem.ram00.INIT_35 = 256'h5CE0307CE05CE04072E076005068E05C0000004E0E124E0000003E0E00313E00,
progmem.ram00.INIT_36 = 256'hBA000096E070B6E09C00BAACE0B000DAA2E096000080E03C92E05E8CE0800000,
progmem.ram00.INIT_37 = 256'hBC00E0D6FAE0EE0000D4E082EAE0EA0012E0E0D40000BAE098D0E0D000DAC6E0,
progmem.ram00.INIT_38 = 256'h000000000000000008E0F02CE02626E00220E0401AE07C14E0080000EEE0F400,
progmem.ram00.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'h003018706C18000000000000000000000000000F00F000000000000000000E1E,
progmem.ram01.INIT_01 = 256'h600000000000003C3C6666663C3C3C42663C3C7E1E103C00003C7E7E3C080000,
progmem.ram01.INIT_02 = 256'h0038384418102004FF0101F0C0FF0000000001041040AA300C00000000000000,
progmem.ram01.INIT_03 = 256'h2808001034083008102000340834280828083810340810300010000038107C00,
progmem.ram01.INIT_04 = 256'h181818546C18000000000000000000000000000F00F028081020003408342808,
progmem.ram01.INIT_05 = 256'h601800000000000C30666666666666666C186060303866001866064066180600,
progmem.ram01.INIT_06 = 256'h1454404420002004FE0302F0C0FF000000FF0104104055181800000000000000,
progmem.ram01.INIT_07 = 256'h0010002858104810281044581058001000104428581000105030000004100000,
progmem.ram01.INIT_08 = 256'h180C1868FE18000000000000000000000000000F00F000102810105810580010,
progmem.ram01.INIT_09 = 256'h66003E3C3E3C000C303C66666066667E781860606038067E18660C7C06380C00,
progmem.ram01.INIT_0A = 256'h286C382820102004FC0704F0C0FF0000000001041040AA181866C6663E3E3CFC,
progmem.ram01.INIT_0B = 256'h383838103838504400002838384438387C7C401000001010281000441C7C0000,
progmem.ram01.INIT_0C = 256'h7E0C00106C18000000000000000000000000000F00F044440044003838580000,
progmem.ram01.INIT_0D = 256'h6C3866666006000C303C7E663C66667E70186E78606C0C00003E0C061C18187E,
progmem.ram01.INIT_0E = 256'h5064447C70101008F80F08F0C0000000FF000104104055066066C666606666D6,
progmem.ram01.INIT_0F = 256'h44444438040478284444104444641010404040101010207C1410104404100038,
progmem.ram01.INIT_10 = 256'h180C002CFE1800000000000000000000000000F0F000444444447C4444643030,
progmem.ram01.INIT_11 = 256'h7818667E603E000C30187E660666666678186660607C187E1806180606183000,
progmem.ram01.INIT_12 = 256'h286C381020101818F01F10F0C0000000000001041040AA181866D6663C6666D6,
progmem.ram01.INIT_13 = 256'h7C7C401C3C3C4410444428444454101070704028282840302810004438100000,
progmem.ram01.INIT_14 = 256'h181800546C0000000000000000000000000000F0F00044444444004444441010,
progmem.ram01.INIT_15 = 256'h6C183E606066000C30186666666E66666C18666030C60000180C186666186000,
progmem.ram01.INIT_16 = 256'h1454047C201007E0E03F20F0C00000FF0000010410405518183ED666063E66C6,
progmem.ram01.INIT_17 = 256'h404044644444641044444444444C101040404444444444085000006400000000,
progmem.ram01.INIT_18 = 256'h0030001C6C1800000000000000000000000000F0F0003C3C4444104444441010,
progmem.ram01.INIT_19 = 256'h663C063C3E3A7E3C3C18423C3C3C3C66663C3C7E1EC618001038183C3C3C0000,
progmem.ram01.INIT_1A = 256'h003838105C100000C07F40F0C0000000000001041040AA300C067C3A7C063CC6,
progmem.ram01.INIT_1B = 256'h3838383C3C3C581038380038384438387C7C387C7C7C38100000005C007C0000,
progmem.ram01.INIT_1C = 256'h00000000000000000000000000000000000000F0F00004043838003838443838,
progmem.ram01.INIT_1D = 256'h00003C0000000000000000000006000000000000000000002000000000000000,
progmem.ram01.INIT_1E = 256'h000000000000000080FF80F0C000FF000000010410405500003C000000060000,
progmem.ram01.INIT_1F = 256'h0000600000008000000000000000000000006044444400380000004000000000,
progmem.ram01.INIT_20 = 256'h34322F2D2A282523201E1B191614110F0C0A0705020038380000000000000000,
progmem.ram01.INIT_21 = 256'h02020202020101010101010101000000000000000046444239373533313C3937,
progmem.ram01.INIT_22 = 256'h0606060606050505050505050504040404040404040303030303030303020202,
progmem.ram01.INIT_23 = 256'h0A0A0A0A0A090909090909090908080808080808080707070707070707060606,
progmem.ram01.INIT_24 = 256'h0E0E0E0E0E0D0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0A0A0A,
progmem.ram01.INIT_25 = 256'h8015010012091300E00900130000120000110913000F0F0F0F0F0F0F0F0E0E0E,
progmem.ram01.INIT_26 = 256'h120841000012091300E009001300001200610000120913000912091E09091109,
progmem.ram01.INIT_27 = 256'h1300091230000009178000120913002E090000110912098015FF001209130009,
progmem.ram01.INIT_28 = 256'h178000120A13002E0A0000110A120A8015FF00120A13000912090A11090A1109,
progmem.ram01.INIT_29 = 256'h090A11000012090A110A0A110A13000A120A0A110A0A110A13000A123000000A,
progmem.ram01.INIT_2A = 256'h0A0013000012000114002B0000120A1300E00A00130000110A13000A3100C041,
progmem.ram01.INIT_2B = 256'h1E0A0A110B80150100120A1300E00A001300001200001400230000120A1300E0,
progmem.ram01.INIT_2C = 256'h0B13000B12090B1100C0110B13000B120A0B11000214C000C0110B13000A120A,
progmem.ram01.INIT_2D = 256'h0B13000B12090B11090B11090B11090B11090B11090B11090B11090B110A0B11,
progmem.ram01.INIT_2E = 256'h0A0B110A0B110A0B110A0B110A0B110A0B110A0B110B1300E00B001300000011,
progmem.ram01.INIT_2F = 256'h14000C170000120B13000B12090B110B0B110B13000B120A0B110A0B110A0B11,
progmem.ram01.INIT_30 = 256'h000C170000120B0C110C13002E0C0000110B0C110C13000B120B0C110B120000,
progmem.ram01.INIT_31 = 256'h0C0C110000110C13000C120C0C1100A108001A0C13000C120C0C110C12000014,
progmem.ram01.INIT_32 = 256'h1A0C13000C120C0C1100A108001A0C13000C120C0C11001B00001A0C13000C12,
progmem.ram01.INIT_33 = 256'hE00C0013FF00120C1300E00C001600B01A0C1300E00CB01B0C0C110C0C1100B0,
progmem.ram01.INIT_34 = 256'h002E0D0000110D13000D00110D00110D00120C0D110D13002E0D0010110D1300,
progmem.ram01.INIT_35 = 256'h0D120D0D110D120D0D110D170D0D110D1300E00D00120D13002E0D0000110D13,
progmem.ram01.INIT_36 = 256'h0D13000D120C0D110D1E0C0D110D170C0D110D13000D120B0D110D0D110D1300,
progmem.ram01.INIT_37 = 256'h0D0E110D0D110D13000D120D0D110D170D0D110D13000D120D0D110D170C0D11,
progmem.ram01.INIT_38 = 256'h00000000000000000E120D0E110B0E110D0E110D0E110B0E110E13000D120D1E,
progmem.ram01.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
