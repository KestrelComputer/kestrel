`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,
	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB00);		// B000-B003 : KIA (B004-BFFF = repeats)
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)};
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h3C1C0C3C180000000C3818660000000000000000000000000000000F0000D600,
progmem.ram00.INIT_01 = 256'h0000080000001800601C06603018007E66C67E7C7C666006667E787C3C200400,
progmem.ram00.INIT_02 = 256'h007C08381038003828100010000000FF8080E0FFFF000000FF02082080361800,
progmem.ram00.INIT_03 = 256'h022810204810201020002810102028083C28102070102010202E281020C03038,
progmem.ram00.INIT_04 = 256'h66301C6624000024186C3E660000000000000000000000000000000F00402808,
progmem.ram00.INIT_05 = 256'h0000180000001818603006601818600666C618666676600666606C6666300C18,
progmem.ram00.INIT_06 = 256'h00F410042874001C001044380000007FC040E0FFFF00000000020820806C1800,
progmem.ram00.INIT_07 = 256'h3C0028103028102810000028082000104C002810482810281058002810201044,
progmem.ram00.INIT_08 = 256'h66603C0666000018306858240000000000000000000000000000000F00400010,
progmem.ram00.INIT_09 = 256'h66663C5E7C5C18007C303E7C0C3C300C3C6C186666766006666066666E181818,
progmem.ram00.INIT_0A = 256'h00F40018106C7C64001038540007E03FE020E0FF000000FF000208208000187E,
progmem.ram00.INIT_0B = 256'h4C38383808000038386C383838380000543838384438387C7C58000000C41044,
progmem.ram00.INIT_0C = 256'h3C7C6C0C6600007E30323C000000000000000000000000000000000F00584444,
progmem.ram00.INIT_0D = 256'h3C66186066661818667C6666003C1818186C187C7C7E60067E78667C6A0C3000,
progmem.ram00.INIT_0E = 256'h007400200074043C000028500018181FF010E0FF00000000000208208000180C,
progmem.ram00.INIT_0F = 256'h5444444438303044441204040424444454444444E4101040408C101010287C38,
progmem.ram00.INIT_10 = 256'h66667E3066001018306C1A0000000000000000000000000000000F0000644444,
progmem.ram00.INIT_11 = 256'h183C1860666618186630666600660C303C381878606E60666660666666181800,
progmem.ram00.INIT_12 = 256'h0014003C006C007C001038540010080FF808E0000000FF000002082080001818,
progmem.ram00.INIT_13 = 256'h644444444410107C7C7E3C3C3C384444544444444410106070F8282828D40800,
progmem.ram00.INIT_14 = 256'h66660C6024181824186C7C0000000000000000000000000000000F0000644444,
progmem.ram00.INIT_15 = 256'h3C3C18607C66181866306666000006606638186C606E606666606C6660300C18,
progmem.ram00.INIT_16 = 256'h00140000006C00000010443800200407FC04E000000000000002082080001830,
progmem.ram00.INIT_17 = 256'h78444444441010404090444444204444644444444810104040884444442C287C,
progmem.ram00.INIT_18 = 256'h3C3C0C7E181810000C3A180000000000000000000000000000000F0000584444,
progmem.ram00.INIT_19 = 256'h66180C6060660C1866303E7C0000007E6610186660667E3C6660787C3C200418,
progmem.ram00.INIT_1A = 256'h08140000003800000010001000200403FE02E00000FF0000000208208000187E,
progmem.ram00.INIT_1B = 256'h8038383838383838386E3C3C3C203838783838387038387C7C8E7C7C7C5C3800,
progmem.ram00.INIT_1C = 256'h00000000000020000000000000000000000000000000000000000F0000403838,
progmem.ram00.INIT_1D = 256'h0000000060000070000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_1E = 256'h10000000000000000000000000200401FF01E000000000000002082080000000,
progmem.ram00.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000444444040800,
progmem.ram00.INIT_20 = 256'h000000000000000000000070009020B040D060F08010A030C050E07000400000,
progmem.ram00.INIT_21 = 256'h0064E06A004C76E07A3A17640000004A3A12023A143A00234A000040E0400000,
progmem.ram00.INIT_22 = 256'hAE3C12063E14AE0000922E3A0041013216809EE09200007EE006423434127E00,
progmem.ram00.INIT_23 = 256'hB000E0003E36A194F2E0E6000000C23A12503A143C00133C123A3CA1C2000000,
progmem.ram00.INIT_24 = 256'hE840E0340000E6E0C430E0C42AE0C424E0C41EE0C418E0C412E0C40CE0C406E0,
progmem.ram00.INIT_25 = 256'h005632503100563812FF38143668E076381756000034E0320113323612013614,
progmem.ram00.INIT_26 = 256'h3041B6000096E09C0058AEE0B20017B0321496000080E06692E03A0030800000,
progmem.ram00.INIT_27 = 256'h00EE2E033014EE0000DAE0B8EAE00600DA0000C6E0B8D6E00200C60000B62E30,
progmem.ram00.INIT_28 = 256'h3014360000262E013014260000001830A118000000FE3031043014F00AE0FE00,
progmem.ram00.INIT_29 = 256'h301476000066E02872E0660000562E043014560000462E023014460000362E02,
progmem.ram00.INIT_2A = 256'h000086E098B8E0360413303812F0A6E03400289CE032003892E0860000762E06,
progmem.ram00.INIT_2B = 256'h1538FEE0F20000BCE042EEE0360413303812F0DCE0340028D2E0320038C8E0BC,
progmem.ram00.INIT_2C = 256'h171A3EE04E0000D815382EE0220000F2E0881EE0F2E01810171A0EE01E0000B0,
progmem.ram00.INIT_2D = 256'h82E05CE0C878E07C0040F0161A68E05C000052E052000022E0BE4EE022E04811,
progmem.ram00.INIT_2E = 256'hB8C0E0080088B6E090E05EACE0B00030F0161A9CE090000086E08600005CE0DC,
progmem.ram00.INIT_2F = 256'h00CEE0DCFAE0C6F4E0CEE092EAE0EE0020F0161ADAE0CE0000C4E0C4000090E0,
progmem.ram00.INIT_30 = 256'h10F0161A3AE02E0000FEE0242AE0F424E02A0000EE152814E02A00F00AE0FE00,
progmem.ram00.INIT_31 = 256'hC880E05EE03076E07A00171A6AE05E00002EE0005AE00054E02EE0D04AE04E00,
progmem.ram00.INIT_32 = 256'h0060BEE0C201171AB2E086ACE0A0000084E0B89CE0019C100130158400005EE0,
progmem.ram00.INIT_33 = 256'hE0CEFEE082F8E0EC0000CC2E30004100142C2C12020042CC0000A0E0C8C8E0A6,
progmem.ram00.INIT_34 = 256'h24482C1732000008E0002C2C41012E71000141FF2A16012C14080000ECE0A204,
progmem.ram00.INIT_35 = 256'h8412692E16700000005C2C12FF2A145C0000004C2C00314C000032E02C002CFF,
progmem.ram00.INIT_36 = 256'h16B8000094E0EEB4E04EAEE00094A8126C2E1694000070E0EE90E05E8AE00070,
progmem.ram00.INIT_37 = 256'hDCE0EEFCE034F6E000DCF0127D2E16DC0000B8E0EED8E00AD2E000B8CC127A2E,
progmem.ram00.INIT_38 = 256'h3A000024E0022E1B000216240000001002122E021310000000E02A0013000000,
progmem.ram00.INIT_39 = 256'h0050E0267AE03C74E0020050E01266E06A00F002165000003AE0404C1E010015,
progmem.ram00.INIT_3A = 256'hBAC0E0DEBAE080B4E0A800007EE084021E7EE0529AE09E00E002163C8AE07E00,
progmem.ram00.INIT_3B = 256'h0000000000D4E0AAF2E0EEECE04EE6E002E0E0D40000A8E0AE0072CCE096C6E0,
progmem.ram00.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'h3C7E7E3C080000003018706C18000000000000000000000000000F00F0000E1E,
progmem.ram01.INIT_01 = 256'h00000000000000600000000000003C3C6666663C3C3C42663C3C7E1E103C0000,
progmem.ram01.INIT_02 = 256'h10000038107C000038384418102004FF0101F0C0FF0000000001041040AA300C,
progmem.ram01.INIT_03 = 256'h2000340834280828080010340830081020003408342808280838103408103000,
progmem.ram01.INIT_04 = 256'h66064066180600181818546C18000000000000000000000000000F00F0280810,
progmem.ram01.INIT_05 = 256'h00000000000000601800000000000C30666666666666666C1860603038660018,
progmem.ram01.INIT_06 = 256'h300000041000001454404420002004FE0302F0C0FF000000FF01041040551818,
progmem.ram01.INIT_07 = 256'h1010581058001000100028581048102810445810580010001044285810001050,
progmem.ram01.INIT_08 = 256'h660C7C06380C00180C1868FE18000000000000000000000000000F00F0001028,
progmem.ram01.INIT_09 = 256'h66C6663E3E3CFC66003E3C3E3C000C303C66666066667E781860606038067E18,
progmem.ram01.INIT_0A = 256'h1000441C7C0000286C382820102004FC0704F0C0FF0000000001041040AA1818,
progmem.ram01.INIT_0B = 256'h44003838580000383838103838504400002838384438387C7C40100000101028,
progmem.ram01.INIT_0C = 256'h3E0C061C18187E7E0C00106C18000000000000000000000000000F00F0444400,
progmem.ram01.INIT_0D = 256'h66C666606666D66C3866666006000C303C7E663C66667E70186E78606C0C0000,
progmem.ram01.INIT_0E = 256'h101044041000385064447C70101008F80F08F0C0000000FF0001041040550660,
progmem.ram01.INIT_0F = 256'h447C444464303044444438040478284444104444641010404040101010207C14,
progmem.ram01.INIT_10 = 256'h06180606183000180C002CFE1800000000000000000000000000F0F000444444,
progmem.ram01.INIT_11 = 256'h66D6663C6666D67818667E603E000C30187E660666666678186660607C187E18,
progmem.ram01.INIT_12 = 256'h10004438100000286C381020101818F01F10F0C0000000000001041040AA1818,
progmem.ram01.INIT_13 = 256'h440044444410107C7C401C3C3C44104444284444541010707040282828403028,
progmem.ram01.INIT_14 = 256'h0C186666186000181800546C0000000000000000000000000000F0F000444444,
progmem.ram01.INIT_15 = 256'h3ED666063E66C66C183E606066000C30186666666E66666C18666030C6000018,
progmem.ram01.INIT_16 = 256'h000064000000001454047C201007E0E03F20F0C00000FF000001041040551818,
progmem.ram01.INIT_17 = 256'h44104444441010404044644444641044444444444C1010404044444444440850,
progmem.ram01.INIT_18 = 256'h38183C3C3C00000030001C6C1800000000000000000000000000F0F0003C3C44,
progmem.ram01.INIT_19 = 256'h067C3A7C063CC6663C063C3E3A7E3C3C18423C3C3C3C66663C3C7E1EC6180010,
progmem.ram01.INIT_1A = 256'h00005C007C0000003838105C100000C07F40F0C0000000000001041040AA300C,
progmem.ram01.INIT_1B = 256'h380038384438383838383C3C3C581038380038384438387C7C387C7C7C381000,
progmem.ram01.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000F0F000040438,
progmem.ram01.INIT_1D = 256'h3C00000006000000003C00000000000000000000060000000000000000000020,
progmem.ram01.INIT_1E = 256'h00004000000000000000000000000080FF80F0C000FF00000001041040550000,
progmem.ram01.INIT_1F = 256'h0000000000000000006000000080000000000000000000000060444444003800,
progmem.ram01.INIT_20 = 256'h00000000000000000000003A3733302C2925221E1B1814110D0A060300383800,
progmem.ram01.INIT_21 = 256'h000812081E080811080812081300E00808130008120800110813000812081300,
progmem.ram01.INIT_22 = 256'h08081300081A081300083108C041000812080811081300081208410808120813,
progmem.ram01.INIT_23 = 256'h08091130080812080811081300E0080813000812080114082B080812081300E0,
progmem.ram01.INIT_24 = 256'h0809110913000812080911080911080911080911080911080911080911080911,
progmem.ram01.INIT_25 = 256'h2E09080011E0090813FF08120909110908120913000912080014080813000812,
progmem.ram01.INIT_26 = 256'h08120913000912091E090911098015FF0812091300091208091108C011091300,
progmem.ram01.INIT_27 = 256'h0009A10008120913000912090911001009130009120909110010091300093108,
progmem.ram01.INIT_28 = 256'h08120A13000AA10008120A13002E0A08120A13002E090841000812090A110913,
progmem.ram01.INIT_29 = 256'h08120A13000A120A0A110A13000A210008120A13000A210008120A13000AA100,
progmem.ram01.INIT_2A = 256'h13000A12090A11080014080813090A1108130A0A1108130A0A110A13000AA100,
progmem.ram01.INIT_2B = 256'h140A0A110A13000A12080A11080014080813090A1108130A0A1108130A0A110A,
progmem.ram01.INIT_2C = 256'h160A0B110B1780FF140A0B110B13000A120A0B110A120B00160A0B110B1780FF,
progmem.ram01.INIT_2D = 256'h0B110B12090B110B170000150A0B110B13000B120B13000B120A0B110B120B00,
progmem.ram01.INIT_2E = 256'h090B1100100B0B110B120B0B110B170000150A0B110B13000B120B13000B1209,
progmem.ram01.INIT_2F = 256'h000B12090B110B0B110B120B0B110B170000150A0B110B13000B120B13000B12,
progmem.ram01.INIT_30 = 256'h0000150A0C110C13000B120B0C110A0C110C1780FF140A0C110C17090C110B13,
progmem.ram01.INIT_31 = 256'h090C110C120C0C110C00160A0C110C13000C120A0C110C0C110C120B0C110C17,
progmem.ram01.INIT_32 = 256'h1E0C0C110C00160A0C110C0C110C13000C12090C11000C170008120C13000C12,
progmem.ram01.INIT_33 = 256'h110C0C11090C110C13000C3108102110440808120010110C13000C12090C110C,
progmem.ram01.INIT_34 = 256'h110D08120D13000D1230080812000D51800014FF08120008120D13000C120C0D,
progmem.ram01.INIT_35 = 256'h0D170008120D1300E00D0813FF08120D13002E0D0800110D13000D12081308FF,
progmem.ram01.INIT_36 = 256'h120D13000D120C0D110D0D11E00D0D170008120D13000D120C0D110D0D11E00D,
progmem.ram01.INIT_37 = 256'h0D120C0D110D0D11E00D0D170008120D13000D120C0D110D0D11E00D0D170008,
progmem.ram01.INIT_38 = 256'h0E13000E12B0081380B01A0E1300E00EB01B08B01A0E13000E120810120E1300,
progmem.ram01.INIT_39 = 256'h000E120E0E110E0E11B01B0E120E0E110E1700B01A0E13000E120E0E1700B01A,
progmem.ram01.INIT_3A = 256'h0D0E110D0E110E0E110E13000E120EB01B0E120E0E110E1700B01A0E0E110E13,
progmem.ram01.INIT_3B = 256'h00000000000E120E0E110C0E110D0E110E0E110E13000E120E1E0D0E110D0E11,
progmem.ram01.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram10.INIT_00 = 256'h531F10326C72734B72666E6961697041747246191032454F534C4D231001C610,
progmem.ram10.INIT_01 = 256'h6475726B61202D657465206D53001001322D652D31322310496F6C462E20656D,
progmem.ram10.INIT_02 = 256'h726F5004102A02107473657520316561742834365374623620554304102A0210,
progmem.ram10.INIT_03 = 256'h20656F686F6F206F645604102A0210293220746562646178284B313A726D6D6D,
progmem.ram10.INIT_04 = 256'h2F5004102A02104B313A726D6D6F645604102A02106C6F736970722065706D69,
progmem.ram10.INIT_05 = 256'h6167722020303002106120726D4D326C72734B00100165617274696461626520,
progmem.ram10.INIT_06 = 256'h07107C2020202064736E20203034021020202020202020207C07107C796F6520,
progmem.ram10.INIT_07 = 256'h02107C2020202020202F2020304202107C18107C07107C18107C07107C18107C,
progmem.ram10.INIT_08 = 256'h736C4D746F4100100120202020202020207C07107C20796F6520656920203043,
progmem.ram10.INIT_09 = 256'h6E7469776D726F706E69616E73722020656E5704102A02106C6E67722832656F,
progmem.ram10.INIT_0A = 256'h6F696F2074652061646F20746C6220656E5704102A02107265206F20746F2069,
progmem.ram10.INIT_0B = 256'h6D722074646565726520747420656E5704102A02106569206169727664616C74,
progmem.ram10.INIT_0C = 256'h682C6F6361656120747420656E5704102A021065616F736B6F62647362686166,
progmem.ram10.INIT_0D = 256'h6B6D6F2067756E6C636663702D696D646570692020656E5704102A02106D6E70,
progmem.ram10.INIT_0E = 256'h102A021029746C652832656F736C4D746F41001001736573646C206E72687520,
progmem.ram10.INIT_0F = 256'h652061646E4304102A0210746C207964346E20746F206E686120696E74695704,
progmem.ram10.INIT_10 = 256'h204904102A02106C766974726473624D5204102A021029746173617374282074,
progmem.ram10.INIT_11 = 256'h5104102A02106D6E7369656E682C6E746569206E6373736C72734B6574656165,
progmem.ram10.INIT_12 = 256'h102D6E74656920756220724D00100165697372687520744C4479726464616B69,
progmem.ram10.INIT_13 = 256'h6C20736C4D6E6C612072206E73206C7274657972652072766E74695704102A02,
progmem.ram10.INIT_14 = 256'h74676E6920737073746E6D35276565706F2704102A0210676C646865206F7261,
progmem.ram10.INIT_15 = 256'h6E67697274207465646E69636472656F5304102A02102D202E3270533230206F,
progmem.ram10.INIT_16 = 256'h65736E6673776B6520646C20695404102A0210656173635274206E6D6F706577,
progmem.ram10.INIT_17 = 256'h746E4304102A0210657563725332656F736C4D0010016875682072746C687520,
progmem.ram10.INIT_18 = 256'h696C4D04102A021064736E206C736D2D207444746F206F423204102A0210736E,
progmem.ram10.INIT_19 = 256'h7475746E206C696C6D736668206F6B61206F207565612074736C61206F74636C,
progmem.ram10.INIT_1A = 256'h2A0210644372767220494D04102A0210736C61727631206C4F04102A0210736F,
progmem.ram10.INIT_1B = 256'h20655504102A021072747272744929432865616761206E6D6F20636861470410,
progmem.ram10.INIT_1C = 256'h204B20697369206C7262747520616772206C4604102A0210727672206366656E,
progmem.ram10.INIT_1D = 256'h654304102A021063657270457465706C764432656F736C4D00100121726D6D66,
progmem.ram10.INIT_1E = 256'h776769692065756920724D04102A0210746565206E6F206C746C3A64636D6F6E,
progmem.ram10.INIT_1F = 256'h6572632C656F6C65696465204104102A021065636A6965652074656520652061,
progmem.ram10.INIT_20 = 256'h2061746E2054454306102A041021746565206E786653554804102A0210746373,
progmem.ram10.INIT_21 = 256'h102A041058206561666E20656C7372414B662073734D06102A04102C54454366,
progmem.ram10.INIT_22 = 256'h102A2C10236769734D2E102A2C106965686961727469707274727274694C4706,
progmem.ram10.INIT_23 = 256'h6E6969696565206E6C532E102A2C10726C6E686E672069727265746F656E462E,
progmem.ram10.INIT_24 = 256'h102A0210746E432063657270457465706C764432656F736C4D001001646F206F,
progmem.ram10.INIT_25 = 256'h642C6D74796569652079643404102A02105352576D6F6E65433A6F736C6E4304,
progmem.ram10.INIT_26 = 256'h656820677276206174655304102A021021726E6F2075206F6673636664656973,
progmem.ram10.INIT_27 = 256'h6F667977206E70206D747468206F25386E6820724D04102A0210612020726F20,
progmem.ram10.INIT_28 = 256'h206F66646E614C736F734C0010016F62746E655304102A021064616265206820,
progmem.ram10.INIT_29 = 256'h7372725304102A0210646465204F2063742072745204102A021067696F205831,
progmem.ram10.INIT_2A = 256'h73526620634C04102A021065612074776562736F206C742070616C6673206C6E,
progmem.ram10.INIT_2B = 256'h74206572664504102A02106575617465656161206F7475696E63736972666B61,
progmem.ram10.INIT_2C = 256'h041072696120746F20744C506D6F6E654306102A041067696D726F7064727475,
progmem.ram10.INIT_2D = 256'h74766E69736D746D5306102A0410657365687520666F7073657465724306102A,
progmem.ram10.INIT_2E = 256'h69634D6E206562747075204E06102A041065656E736F74646F206965706F2076,
progmem.ram10.INIT_2F = 256'h29276F2867696F205831206F66646E614C736F734C0010016875682068724665,
progmem.ram10.INIT_30 = 256'h6C4D06102A0410646465206C74727065206F7475746E206C696C4D04102A0210,
progmem.ram10.INIT_31 = 256'h6D74622C734606102A04106C6120756B6F20676F682072746478667920656C69,
progmem.ram10.INIT_32 = 256'h021029276F2867696F205831206F66646E614C736F734C00100179677520726D,
progmem.ram10.INIT_33 = 256'h206561206C634104102A021065656E7965616573646E6963727369524A04102A,
progmem.ram10.INIT_34 = 256'h107C202064416E75657C04107C4F204F204920497C04102E726D6D6620657920,
progmem.ram10.INIT_35 = 256'h537C537C041032796E206561207369524A04102A02107C207365644172757C04,
progmem.ram10.INIT_36 = 256'h614C736F734C0010014D5266204B2E2074656E20765304102A02107C72642062,
progmem.ram10.INIT_37 = 256'h656165736465616F7368614604102A021029276F2867696F205831206F66646E,
progmem.ram10.INIT_38 = 256'h2065776473206C4F06102A04104F206F42327373206E4606102A041065656E79,
progmem.ram10.INIT_39 = 256'h676D204B2068206F4235336561206C6F2020746D74654904102A021067696E72,
progmem.ram10.INIT_3A = 256'h6C3A644504102A02106569737472663A6D4804102A02106F7467764E0010012E,
progmem.ram10.INIT_3B = 256'h646C206E6B4D001001756965703A555004102A0210786E3A445004102A021073,
progmem.ram10.INIT_3C = 256'h656973732E732D646C20746F672404102A021029276F2832656F736C4D726673,
progmem.ram10.INIT_3D = 256'h726F5004102A02104549786969207469736C7372657370744304102A0210732E,
progmem.ram10.INIT_3E = 256'h5104102A02106E4604102A02106F00100174652068206F20706864612C47466D,
progmem.ram10.INIT_3F = 256'h00000000000000000000000000A0F084B08ED2260A4CD6A49830566206014126;

defparam
progmem.ram11.INIT_00 = 256'h61120AE52D657465206F206F74636C702073691F08FF2D4E5445490B07000F00,
progmem.ram11.INIT_01 = 256'h7F6E6F676342326C72734B656F190000BF32705332300B0B4920766120416C75,
progmem.ram11.INIT_02 = 256'h6167722703200203296572707336726D655320583120692D313A502602200202,
progmem.ram11.INIT_03 = 256'h622C6D72636E4D3A65692A04200204844B336F206C616E7045203620796F6520,
progmem.ram11.INIT_04 = 256'h32531706200206FC3620796F652065691105200205796E206368616764706174,
progmem.ram11.INIT_05 = 256'h6D726F507C30301703704D796F65202D657465140000F06366656E20726F796B,
progmem.ram11.INIT_06 = 256'h0106FF20202020206575557C303017057C20202020202020201204EE20726D6D,
progmem.ram11.INIT_07 = 256'h170AFF2020202020204F497C303017092F0108E50108FF0107FF01072F0106F3,
progmem.ram11.INIT_08 = 256'h7465692075621C00007C2020202020202020120BE52020726D4D6F64567C3030,
progmem.ram11.INIT_09 = 256'h2065747220616772206F7474656570616474613802200202296169696F202D6E,
progmem.ram11.INIT_0A = 256'h6E7A72682C787477722074796969616474613A0320020373617972666872466E,
progmem.ram11.INIT_0B = 256'h206F66616120766974726F20696474613904200204736E6C6C637465206E2061,
progmem.ram11.INIT_0C = 256'h69206C6F202076686F206964746122052002050367727420636C2065612D736C,
progmem.ram11.INIT_0D = 256'h656120746561676120696965736E616F206C6D73616474614606200206656120,
progmem.ram11.INIT_0E = 256'h022002020079696172202D6E7465692075621B000079612065697367696F7461,
progmem.ram11.INIT_0F = 256'h7874777220611F03200203FF616673612020696872466569634D6E2065747227,
progmem.ram11.INIT_10 = 256'h627438052002052E616572652065612D4F1404200204F82E727420202749202E,
progmem.ram11.INIT_11 = 256'h7524062002066561207420636520656F736C6D646F6520276574652068206D63,
progmem.ram11.INIT_12 = 256'h0232656F736C4D746F61656F16000073646C206F74616F2053207469206E2063,
progmem.ram11.INIT_13 = 256'h6543276C69206172482E446769757965696E206C616E7965206574724A022002,
progmem.ram11.INIT_14 = 256'h206869646D746120657569202064746C6D433803200203796F6F6F746D6D6F6E,
progmem.ram11.INIT_15 = 256'h65206E7461736F2075206F7475652070633B04200204293A20322D652D31326E,
progmem.ram11.INIT_16 = 256'h64686969206120636465697373683005200205DF63706B6120617465796C6D20,
progmem.ram11.INIT_17 = 256'h61736F09022002020872747574202D6E7465691500002E676F742C656120636D,
progmem.ram11.INIT_18 = 256'h70747549042002042E65757579746F202D6161206E4666204B2203200203D774,
progmem.ram11.INIT_19 = 256'h6963727369797074752F7469736620636C726670206B6D6F206562746E696169,
progmem.ram11.INIT_1A = 256'h200207656F206569444147100620020621656269612031796E1205200205FF6E,
progmem.ram11.INIT_1B = 256'h497273150820020895656570656E204C472067756E4C64616D43736970722B07,
progmem.ram11.INIT_1C = 256'h6F42346E20746679656120736A6D726F706C752F0A20020A0B65694465617274,
progmem.ram11.INIT_1D = 256'h616C2402200202656E696578206E6D6F6565202D6E746569220000A2796F6520,
progmem.ram11.INIT_1E = 256'h68206E786673746E6D65653203200203736366646F207465746920656F206F72,
progmem.ram11.INIT_1F = 256'h726E6F20646D6F206E6C61647320042002046474656E20727773636664776674,
progmem.ram11.INIT_20 = 256'h6F646573694541521906200206FC7363666467696920524F15052002052E7520,
progmem.ram11.INIT_21 = 256'h082002080055796B6C2069647475652049206F6575692307200207F645415220,
progmem.ram11.INIT_22 = 256'h072002072C206E73690A0620020663746D747220656E6F20656570656E204322,
progmem.ram11.INIT_23 = 256'h206F746E6664727465691C08200208F76564612044506E206F7220737063651F,
progmem.ram11.INIT_24 = 256'h0220020229276F28656E696578206E6D6F6565202D6E7465692A000073727766,
progmem.ram11.INIT_25 = 256'h652065692072766C6473612037032002032E4B4F206F72616C206E6975636F1C,
progmem.ram11.INIT_26 = 256'h657274656165616E206E702204200204FF7365726374636D7220746565207470,
progmem.ram11.INIT_27 = 256'h6D722061617465736569206174662030206174656F3705200205796461737568,
progmem.ram11.INIT_28 = 256'h536D7220657265206E73652100006B6F656F20650C0620020624726F796B6574,
progmem.ram11.INIT_29 = 256'h6969707531032002032E65656E544E6B61736E75651802200202DE6E64433436,
progmem.ram11.INIT_2A = 256'h742D206F6B613504200204FF72636869206C6973706C69737370207565757967,
progmem.ram11.INIT_2B = 256'h727364636F6E1F05200205C673622F6E6D676E6D6E69616E746F2064626F2063,
progmem.ram11.INIT_2C = 256'h0207646573656872466F2044206F72616C1D06200206996E6D61677220657563,
progmem.ram11.INIT_2D = 256'h69616F6E206569656F300820020872696120636D736F7220736E63726F1E0720,
progmem.ram11.INIT_2E = 256'h6E68612069736C61206D6A6F2709200209646465206E69696E637478206F6C65,
progmem.ram11.INIT_2F = 256'hF7746E43206E64433436536D7220657265206E736529000000676F742C746F20,
progmem.ram11.INIT_30 = 256'h74752E032002030065656E7965616573646E6963727369797074752702200202,
progmem.ram11.INIT_31 = 256'h6520752074611704200204656274702D6F6C687572746D652065692062736970,
progmem.ram11.INIT_32 = 256'h020200746E43206E64433436536D7220657265206E736529000000726E68796F,
progmem.ram11.INIT_33 = 256'h36736B746C61201F03200203646465206C74727065206F7475746E2053220220,
progmem.ram11.INIT_34 = 256'h06002020726420727452110500504E2047544C544C110400796F65206F737462,
progmem.ram11.INIT_35 = 256'h7520524A11082E206C6F736B746E6E2053160720020700202073726420625311,
progmem.ram11.INIT_36 = 256'h7265206E7365290000004F206F4235312E732061656119092002090020644172,
progmem.ram11.INIT_37 = 256'h6C747270652067727420736C200220020200746E43206E64433436536D722065,
progmem.ram11.INIT_38 = 256'h706E68206575796E17042002044D5266204B206575746F140320020364646520,
progmem.ram11.INIT_39 = 256'h6561694234657466204B2E2076736475634965616973202F05200205006E7469,
progmem.ram11.INIT_3A = 256'h6120206E0A032002032E646C20736920656F12022002026E696169610A000000,
progmem.ram11.INIT_3B = 256'h656953676961250000736F76722070670E052002057465206E670A0420020474,
progmem.ram11.INIT_3C = 256'h73646C20666D61656973687266201F0220020200746E63202D6E746569206F20,
progmem.ram11.INIT_3D = 256'h61677224042002040044206E6C586F6E207475652074612F7521032002030066,
progmem.ram11.INIT_3E = 256'h2005032002032E6904022002026B0200002E736265747266656F206E20415020,
progmem.ram11.INIT_3F = 256'h000000000000000000000000000F0E0E0D0C0B0A090705040302010000000020;

endmodule
