`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,

	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO,
	
	// SD Card Interface
	output			N2_SD_CLK_O,
	output			N2_SD_MOSI_O,
	output			N2_SD_CS_O,
	output			N2_SD_LED_O,

	input				N2_SD_MISO_I,
	input				N2_SD_WP_I,
	input				N2_SD_CD_I
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				gpia_ack_o;
	wire	[15:0]	gpia_dat_o;
	wire				gpia_stb_i;
	wire	[15:0]	gpia_port_o;

	assign N2_SD_CLK_O	= gpia_port_o[3];
	assign N2_SD_MOSI_O	= gpia_port_o[2];
	assign N2_SD_CS_O		= gpia_port_o[1];
	assign N2_SD_LED_O	= gpia_port_o[0];

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB00);		// B000-B003 : KIA
	assign gpia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB01);		// B010-B013 : GPIA 
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i & ~gpia_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	wire	[15:0]	gpia_mask			= {16{gpia_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)} | (gpia_mask & gpia_dat_o);
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | (gpia_stb_i & gpia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	GPIA gpia(
		.RST_I(N2_BTN0_I),
		.CLK_I(mgia_25mhz_o),
		.ADR_I(cpu_adr_o[1]),
		.CYC_I(cpu_cyc_o),
		.STB_I(gpia_stb_i),
		.WE_I(cpu_we_o),
		.DAT_I(cpu_dat_o),
		.DAT_O(gpia_dat_o),
		.ACK_O(gpia_ack_o),
		.PORT_I({13'h0000, N2_SD_MISO_I, N2_SD_WP_I, N2_SD_CD_I}),
		.PORT_O(gpia_port_o)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h03ABABAB03FF0000000000000000000000000000000000000000B600D8001600,
progmem.ram00.INIT_01 = 256'h0D1015740000FF6BCB8BCB6BF303030303ABABAB03FFFF0B0B0B0B0BF3030303,
progmem.ram00.INIT_02 = 256'h15B8000000A41212F71215A4000094E00C101594000084E003101584000074E0,
progmem.ram00.INIT_03 = 256'hBA00E0F4000000E01212081216E0000000CC1212FD1215CC000000B81212FB12,
progmem.ram00.INIT_04 = 256'h1438000028E0041015280000000E1212021216CE1AE00E000000F41212041216,
progmem.ram00.INIT_05 = 256'h6AE03A7CE01403306A000054E03A66E014E83054000038E03E501E141412FF14,
progmem.ram00.INIT_06 = 256'h802415B4000096E0BAB0E096E0F6A6E0AA0096000080E0E292E06C8CE0800000,
progmem.ram00.INIT_07 = 256'hE0B6FEE0B6F8E0B6F2E0B6ECE0E0000000B424B124241A82D2E082CCE098C6E0,
progmem.ram00.INIT_08 = 256'h1AE0E23CE0242E1BE230E02400012E4A1A0000E0E0B616E0B610E0B60AE0B604,
progmem.ram00.INIT_09 = 256'h7A000040E0E276E0241F1B1C6AE02E20131C5EE02E2213E252E0241E1B400000,
progmem.ram00.INIT_0A = 256'h3196161E16FF2482B2E082ACE0BE002AA2E0C816179000007AE0E28CE024FFB0,
progmem.ram00.INIT_0B = 256'h4200E0F40000D2E092F0E0F6EAE0160000300031D20000009030013100903000,
progmem.ram00.INIT_0C = 256'h00002CE00126152C0000001801120C24E0180000000A30120A0000F4E0D406E0,
progmem.ram00.INIT_0D = 256'h74261274000000600112526CE060000050E0042615500000003C01122E48E03C,
progmem.ram00.INIT_0E = 256'h82C0E082BAE025011B25B41A2AA8E025B025251A92000082E000281582000000,
progmem.ram00.INIT_0F = 256'h9400E094FAE094F4E094EEE094E8E094E2E094DCE094D6E02500B0C4000092E0,
progmem.ram00.INIT_10 = 256'h1AE02C251BC636E000012C2511C626E01A000004E026251BC610E0040000C4E0,
progmem.ram00.INIT_11 = 256'h82E000627C127C2615066EE062000040E02A2C131C58E0282C131C4CE0400000,
progmem.ram00.INIT_12 = 256'h180141181A31011A211A2512C6A8E0CE321796000086E06492E086000062E042,
progmem.ram00.INIT_13 = 256'hE80212FF2516C6F4E0E80000D2E098E4E0320030D2000096E0009C3231FF3221,
progmem.ram00.INIT_14 = 256'h002C40127638E02C00000AE0C628E0C622E0D41CE0EA16E00A0000E8E0EE0000,
progmem.ram00.INIT_15 = 256'hE01F95B04C78E01E40B0CE6CE0600000004A2212002000314A00002CE00C46E0,
progmem.ram00.INIT_16 = 256'hC2E04CBCE01E41B0CEB0E0A4000060E07CA0E0109AE00694E094001A8AE0F684,
progmem.ram00.INIT_17 = 256'h8720114CFAE01E48B0CEEEE0E20000A4E07CDEE010D8E006D2E0D2001AC8E0F6,
progmem.ram00.INIT_18 = 256'h11001E50B1CE36E02A0000E2E07C26E01020E0881AE01A001A10E0F60AE0001F,
progmem.ram00.INIT_19 = 256'h1E51B0CE7AE06E00002AE07C6AE01064E0065EE05E001A54E0F64EE000220020,
progmem.ram00.INIT_1A = 256'hE0B800006EE07CB4E010AEE02EA8E006A2E0A8001A98E0F692E0201C134C86E0,
progmem.ram00.INIT_1B = 256'h02E0F60000B8E07CF2E010ECE006E6E0E6001ADCE0F6D6E04CD0E01E77B0CEC4,
progmem.ram00.INIT_1C = 256'hF640E00020002211F830E01E69B0CE24E0BA1EE0120000F6002E00F6000C1196,
progmem.ram00.INIT_1D = 256'hE0F67EE04C78E01E7AB0CE6CE060000012E07C5CE01056E00650E050001A46E0,
progmem.ram00.INIT_1E = 256'hC2E07CBCE07CB6E07CB0E07CAAE09E000060E07C9AE01094E0648EE08E001A84,
progmem.ram00.INIT_1F = 256'h02E010FCE0F6F6E0A6F0E0E400009EE07CE0E07CDAE07CD4E07CCEE07CC8E07C,
progmem.ram00.INIT_20 = 256'h7040E01C12137034E0001C001811001A003116000000060E0131060000E4E0A0,
progmem.ram00.INIT_21 = 256'hE0087EE07E007674E044E0086AE06E000C60E02C5AE044E0540E1744000016E0,
progmem.ram00.INIT_22 = 256'h00A8E084BAE0100430A800000092121201100831920000008212003182000044,
progmem.ram00.INIT_23 = 256'h02E0060084F8E0BEE008EEE0F20076E4E0BEE008DAE0DE000CD0E062CAE0BE00,
progmem.ram00.INIT_24 = 256'h0010E0C03AE010E08430E034008626E010E0200E17100000BEE0AA0CE0BEE094,
progmem.ram00.INIT_25 = 256'hE0087EE082000C74E0406EE06200003EE0A65EE03EE01454E058000110163E00,
progmem.ram00.INIT_26 = 256'h86E008BCE0C00076B2E0D20052A8E064A2E0569CE086E0960E1786000062E062,
progmem.ram00.INIT_27 = 256'hE0020E17F2000086E008EEE0EE0076E4E08CDE1E2ED8E08CE01001D21186C6E0,
progmem.ram00.INIT_28 = 256'h4611523CE0300000F2E0082CE02C005222E0F2E00818E01C000C0EE06208E0F2,
progmem.ram00.INIT_29 = 256'h1012327CE04CE00872E076000C68E0E462E04CE05C0E174C0000300C2E003003,
progmem.ram00.INIT_2A = 256'h31B8000084E008B4E0B4003EAAE084E008A0E0A4000C96E06290E0840000004C,
progmem.ram00.INIT_2B = 256'hE046FEE012F8E088F2E0F4ECE04EE6E086E0E002002AD6E0E6D0E00E00001000,
progmem.ram00.INIT_2C = 256'h0E40E01C00302E00000CE0121C1E021C141C00232A1C170C0000B8E00808E0B8,
progmem.ram00.INIT_2D = 256'h4680E0467AE04674E068000000441C12501C141A02131A121C1A214400002EE0,
progmem.ram00.INIT_2E = 256'hE08CBEE01C3630AC00008AE06AA8E06AA2E06A9CE06A96E08A000068E04686E0,
progmem.ram00.INIT_2F = 256'h1212011216D8F6E0EA000000D61212FE1215D6000000C20112011015C20000AC,
progmem.ram00.INIT_30 = 256'hAE40E01A34303034E0D82EE022000004E00A00041AE01A00C410E004000000EA,
progmem.ram00.INIT_31 = 256'h0017188E12C476E01870E06400004AE00000305CE0D856E04A000022E00646E0,
progmem.ram00.INIT_32 = 256'hD8C0E0B4000098E024B0E09EAA1EC4A4E098000064E02494E04C8EE00888E088,
progmem.ram00.INIT_33 = 256'hE004000E0A12C4F4E0BAEEE030E8E0ECE2E0D60000B4E09AD2E0AECCE01A5430,
progmem.ram00.INIT_34 = 256'h00000014E02436E00430E03000C426E03020E0140000D6E02410E0660AE00804,
progmem.ram00.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'hC8CA6232180F000000000000FE000000000000000000000000000C1E0C1E0D1E,
progmem.ram01.INIT_01 = 256'h000012001300FFD6D3D1D3D6CFC0C0C8C8CA6232180FFFD0D0D0D0D0CFC0C0C8,
progmem.ram01.INIT_02 = 256'h12001300E000B013FFB012001300001200001200130000120000120013000012,
progmem.ram01.INIT_03 = 256'h000111001300E000B01300B012001300E000B013FFB012001300E000B013FFB0,
progmem.ram01.INIT_04 = 256'h12011300011200B012011300E001B01300B012000111011300E000B01300B012,
progmem.ram01.INIT_05 = 256'h011201011100001101130001120101110003110113000112010117000013FF00,
progmem.ram01.INIT_06 = 256'h00001A0113000112000111011200011101170113000112000111010111011300,
progmem.ram01.INIT_07 = 256'h110101110101110101110101110113002E01004100001A010111010111010111,
progmem.ram01.INIT_08 = 256'h021201021100001A010211001B00001102130001120102110102110102110102,
progmem.ram01.INIT_09 = 256'h021300021201021100001A02021100001202021100001201021100001A021300,
progmem.ram01.INIT_0A = 256'h1102001300FF1101021101021102170102110200120213000212010211000011,
progmem.ram01.INIT_0B = 256'h02031102130002120202110002110013200000110213002E020000112E020000,
progmem.ram01.INIT_0C = 256'h1300031200001A031300E0030016030311031300E00300120313000212020311,
progmem.ram01.INIT_0D = 256'h03001A031300E0030016030311031300031200001A031300E003001603031103,
progmem.ram01.INIT_0E = 256'h010311010311000016000317010311004100001A0313000312400012031300E0,
progmem.ram01.INIT_0F = 256'h0304110303110303110303110303110303110303110303110000110313000312,
progmem.ram01.INIT_10 = 256'h041200001A0304114B0000001A030411041300041200001A0304110413000312,
progmem.ram01.INIT_11 = 256'h0411E004041700001A0404110413000412000012040411000012040411041300,
progmem.ram01.INIT_12 = 256'h0000210000410000B100001A0304110400120413000412040411041300041204,
progmem.ram01.INIT_13 = 256'h04051700001A03041104130004120404110002110413000412E0040041FF0031,
progmem.ram01.INIT_14 = 256'hE005051703051105130005120305110305110405110405110513000412041EE0,
progmem.ram01.INIT_15 = 256'h11000011050511000011000511051300E0050013000000110513000512050511,
progmem.ram01.INIT_16 = 256'h0511050511000011000511051300051202051101051104051105170305110205,
progmem.ram01.INIT_17 = 256'h0000130505110000110005110513000512020511010511040511051703051102,
progmem.ram01.INIT_18 = 256'h130200001100061106130005120206110106110406110617030611020611B000,
progmem.ram01.INIT_19 = 256'h0000110006110613000612020611010611040611061703061102061130000000,
progmem.ram01.INIT_1A = 256'h1106130006120206110106110506110406110617030611020611000012050611,
progmem.ram01.INIT_1B = 256'h0711061300061202061101061104061106170306110206110506110000110006,
progmem.ram01.INIT_1C = 256'h02071130000000130607110000110007110607110713000600112E0640071700,
progmem.ram01.INIT_1D = 256'h1102071105071100001100071107130007120207110107110407110717030711,
progmem.ram01.INIT_1E = 256'h0711020711020711020711020711071300071202071101071104071107170307,
progmem.ram01.INIT_1F = 256'h0811010711000711000711071300071202071102071102071102071102071102,
progmem.ram01.INIT_20 = 256'h060811000012060811300000001300003C110813002E08000011081300071207,
progmem.ram01.INIT_21 = 256'h1208081108170308110812080811081703081106081108120800120813000812,
progmem.ram01.INIT_22 = 256'h000812080811000011081300E0080013000000110813002E0800021108130008,
progmem.ram01.INIT_23 = 256'h0911091703081108120808110817030811081208081108170308110708110813,
progmem.ram01.INIT_24 = 256'h0009120809110912080911091700091109120900120913000812080911081208,
progmem.ram01.INIT_25 = 256'h1208091109170309110909110913000912050911091207091109170000120913,
progmem.ram01.INIT_26 = 256'h0912080911091700091109170309110909110109110912090012091300091209,
progmem.ram01.INIT_27 = 256'h120A001209130009120809110917030911090917030911093100000917000911,
progmem.ram01.INIT_28 = 256'h0A17030A110A13000912080A110A17030A110912080A110A17030A11070A1109,
progmem.ram01.INIT_29 = 256'h00130A0A110A12080A110A17030A11050A110A120A00120A13000A00112E0A00,
progmem.ram01.INIT_2A = 256'h110A13000A12080A110A17030A110A12080A110A17030A11050A110A1300E00A,
progmem.ram01.INIT_2B = 256'h12080A11090A11090A11090A110A0A110A0A110B17010A11070A110013000000,
progmem.ram01.INIT_2C = 256'h0B0B1100C0110B13000B120B00130000120000110B00120B13000A12080B110A,
progmem.ram01.INIT_2D = 256'h0B0B110B0B110B0B110B1300E00B001300001200001400230000120B13000B12,
progmem.ram01.INIT_2E = 256'h120B0B1100D3110B13000B120B0B110B0B110B0B110B0B110B13000B120B0B11,
progmem.ram01.INIT_2F = 256'hB01300B0120B0B110B1300E00BB013FFB0120B1300E00B001600B0120B13000B,
progmem.ram01.INIT_30 = 256'h0B0C110000110B0C110B0C110C13000C120C1E000C110C170B0C110C1300E00B,
progmem.ram01.INIT_31 = 256'h0416000C170B0C11080C110C13000C123C1E0B0C110B0C110C13000C120C0C11,
progmem.ram01.INIT_32 = 256'h0B0C110C13000C120C0C110C0C170B0C110C13000C120C0C110C0C11000C110C,
progmem.ram01.INIT_33 = 256'h110D17000D170B0C110A0C110B0C110B0C110C13000C120C0C110B0C11000011,
progmem.ram01.INIT_34 = 256'h0000000D120C0D11000D110D170B0D110B0D110D13000C120C0D110C0D11000D,
progmem.ram01.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
