`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,

	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO,
	
	// SD Card Interface
	output			N2_SD_CLK_O,
	output			N2_SD_MOSI_O,
	output			N2_SD_CS_O,
	output			N2_SD_LED_O,

	input				N2_SD_MISO_I,
	input				N2_SD_WP_I,
	input				N2_SD_CD_I
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				gpia_ack_o;
	wire	[15:0]	gpia_dat_o;
	wire				gpia_stb_i;
	wire	[15:0]	gpia_port_o;

	assign N2_SD_CLK_O	= gpia_port_o[3];
	assign N2_SD_MOSI_O	= gpia_port_o[2];
	assign N2_SD_CS_O		= gpia_port_o[1];
	assign N2_SD_LED_O	= gpia_port_o[0];

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB00);		// B000-B003 : KIA
	assign gpia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB01);		// B010-B013 : GPIA 
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i & ~gpia_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	wire	[15:0]	gpia_mask			= {16{gpia_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)} | (gpia_mask & gpia_dat_o);
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | (gpia_stb_i & gpia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	GPIA gpia(
		.RST_I(N2_BTN0_I),
		.CLK_I(mgia_25mhz_o),
		.ADR_I(cpu_adr_o[1]),
		.CYC_I(cpu_cyc_o),
		.STB_I(gpia_stb_i),
		.WE_I(cpu_we_o),
		.DAT_I(cpu_dat_o),
		.DAT_O(gpia_dat_o),
		.ACK_O(gpia_ack_o),
		.PORT_I({13'h0000, N2_SD_MISO_I, N2_SD_WP_I, N2_SD_CD_I}),
		.PORT_O(gpia_port_o)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h0303ABABAB03FF0000000000000000000000000000000000000066008800CC00,
progmem.ram00.INIT_01 = 256'hE00D1015720000FF6BCB8BCB6BF303030303ABABAB03FFFF0B0B0B0B0BF30303,
progmem.ram00.INIT_02 = 256'h12F71215B2000000A218FF31A2000092E00C101592000082E003101582000072,
progmem.ram00.INIT_03 = 256'hEE1212081216EE000000DA1212FD1215DA000000C61212FB1215C6000000B212,
progmem.ram00.INIT_04 = 256'hE00410153200001C2E121261DC28E01C000000021212041216C80EE002000000,
progmem.ram00.INIT_05 = 256'h1464307400005EE04470E014E8305E000042E0485A1E141412FF141442000032,
progmem.ram00.INIT_06 = 256'h00A0E0C8BAE0A0E004B0E0B400A000008AE0F09CE07696E08A000074E04486E0,
progmem.ram00.INIT_07 = 256'h02E0C0FCE0C0F6E0EA000000BE24B124241A8CDCE08CD6E0A2D0E0802415BE00,
progmem.ram00.INIT_08 = 256'h242E1BEC3AE02400012E4A240000EAE0C020E0C01AE0C014E0C00EE0C008E0C0,
progmem.ram00.INIT_09 = 256'hEC80E0241F1B2674E02E20132668E02E2213EC5CE0241E1B4A000024E0EC46E0,
progmem.ram00.INIT_0A = 256'hFF248CBCE08CB6E0C80034ACE0D216179A000084E0EC96E024FFB08400004AE0,
progmem.ram00.INIT_0B = 256'hE0F80000DCE09CF4E004EEE0160030DC0000009A300131009A300031A0161E16,
progmem.ram00.INIT_0C = 256'h25B025251A300000001C01121028E01C0000000E30120E0000F8E0DE0AE04C04,
progmem.ram00.INIT_0D = 256'h3280E0327AE03274E02500B062000030E08C5EE08C58E025011B25521A3446E0,
progmem.ram00.INIT_0E = 256'h32C0E032BAE02500B0A8000062E026251B329EE03298E03292E0328CE03286E0,
progmem.ram00.INIT_0F = 256'hE000012C2511AAF4E0E80000A8E032E4E032DEE032D8E032D2E032CCE032C6E0,
progmem.ram00.INIT_10 = 256'h2615643CE03000000EE02A2C13EA26E0282C13EA1AE00E0000E8E02C251BAA04,
progmem.ram00.INIT_11 = 256'h7A0000006422120020003164000054E03260E054000030E01050E000304A127C,
progmem.ram00.INIT_12 = 256'h007AE086BAE01EB4E064AEE0AE001EA4E0FA9EE01F95B06692E01E40B0DC86E0,
progmem.ram00.INIT_13 = 256'h0000BEE086F8E01EF2E064ECE0EC001EE2E0FADCE066D6E01E41B0DCCAE0BE00,
progmem.ram00.INIT_14 = 256'h00FCE0863AE01E34E0562EE02E001E24E0FA1EE020006614E01E48B0DC08E0FC,
progmem.ram00.INIT_15 = 256'hE0867EE01E78E06472E072001E68E0FA62E00022002011001E50B1DC4AE03E00,
progmem.ram00.INIT_16 = 256'h82E086BCE01EB6E064B0E0B0001EA6E0FAA0E0669AE01E77B0DC8EE08200003E,
progmem.ram00.INIT_17 = 256'h002211C2FAE01E69B0DCEEE084E8E0DC0000C0002E00C000D61194CCE0C00000,
progmem.ram00.INIT_18 = 256'h42E01E7AB0DC36E02A0000DCE08626E01E20E0641AE01A001E10E0FA0AE00020,
progmem.ram00.INIT_19 = 256'hE078000068E00126156800002AE08664E01E5EE03258E058001E4EE0FA48E066,
progmem.ram00.INIT_1A = 256'h0000B02612B00000009C01128EA8E09C00008CE00426158C0000007801126A84,
progmem.ram00.INIT_1B = 256'hE08CFEE08CF8E08CF2E08CECE08CE6E08CE0E08CDAE0CE0000BEE0002815BE00,
progmem.ram00.INIT_1C = 256'hE0D03EE0D038E0D032E0D02CE0D026E0D020E0140000CEE08C10E08C0AE08C04,
progmem.ram00.INIT_1D = 256'h00700E01317000004EE0166CE01E66E00460E0B45AE04E000014E0D04AE0D044,
progmem.ram00.INIT_1E = 256'h72C0E0C600B2B6E000800E013172A6E0B000109CE04096E080E0900E17800000,
progmem.ram00.INIT_1F = 256'h02E0100430F0000000DA121201100831DA000000CA120031CA000080E00E0130,
progmem.ram00.INIT_20 = 256'h0131723CE04600B232E000060E01317222E02C001018E02C12E0060000F0E0CC,
progmem.ram00.INIT_21 = 256'hE08800847AE064E0740E1764000006E0F260E006E0DC56E05A00C04CE000060E,
progmem.ram00.INIT_22 = 256'hC2E0B6000092E0C0B2E092E0DEA8E0AC0001101692000064E0088EE064E0CC84,
progmem.ram00.INIT_23 = 256'h02E0B8FCE060F6E0E0E0F00E17E00000B6E000B60E013172D2E0DC0010C8E094,
progmem.ram00.INIT_24 = 256'h100144118438E000E00EA1317228E03200741EE000E00EF131180C171044128E,
progmem.ram00.INIT_25 = 256'h2C80E06AE07A0E176A0000E0E00E01307260E06600B256E0E6501E6A4AE0E6E0,
progmem.ram00.INIT_26 = 256'h8EC0E0B400006AE00E013072AAE0B0008EA0E0006A0E01317290E09A001086E0,
progmem.ram00.INIT_27 = 256'h00D00E013172F6E0000010ECE0FEE6E0D0E0E00E17D00000B40C2E00B403CA11,
progmem.ram00.INIT_28 = 256'hE04A007A3AE0000E0E0131722AE034001020E07C1AE00E000000D01012B606E0,
progmem.ram00.INIT_29 = 256'h82E0D27CE01076E09800346CE05066E00E00001000314E00000EE00E01307244,
progmem.ram00.INIT_2A = 256'h021C141C0023C61C17A80000004E0EFF31729EE04EE08294E0668EE0E288E06C,
progmem.ram00.INIT_2B = 256'hDE1C12501C141A02131A121C1A21DE0000CAE0AADAE01C00CA0000A8E0AE1C1E,
progmem.ram00.INIT_2C = 256'h42E0043CE00436E00430E024000002E0E020E0E01AE0E014E0E00EE002000000,
progmem.ram00.INIT_2D = 256'h1212FE1215700000005C01120110155C000046E02658E01C363046000024E004,
progmem.ram00.INIT_2E = 256'h00009EE0A40004B4E0B4005EAAE09E0000008412120112167290E08400000070,
progmem.ram00.INIT_2F = 256'hE0F80000DEE00000CCF0E072EAE0DE0000BCE0A0DAE048D4E01A323072C8E0BC,
progmem.ram00.INIT_30 = 256'h125E3EE0320000F8E0BE2EE0E028E00822E00EAA302200171828125E0AE0A404,
progmem.ram00.INIT_31 = 256'h82E0487CE01A52307270E064000032E0BE60E0380052FF1B26021A26001A0E5A,
progmem.ram00.INIT_32 = 256'hFAC0E008BAE0000ECCBA110EC0125EA4E0509EE0CC98E08692E086000064E034,
progmem.ram00.INIT_33 = 256'h0000000000000000CAE0BEECE004E6E0E6005EDCE0CCD6E0CA000086E0BEC6E0,
progmem.ram00.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'hC8C8CA6232180F000000000095000000000000000000000000000C1E0C1E0C1E,
progmem.ram01.INIT_01 = 256'h12000012001300FFD6D3D1D3D6CFC0C0C8C8CA6232180FFFD0D0D0D0D0CFC0C0,
progmem.ram01.INIT_02 = 256'h13FFB0120013002E000003110013000012000012001300001200001200130000,
progmem.ram01.INIT_03 = 256'h00B01300B012001300E000B013FFB012001300E000B013FFB012001300E000B0,
progmem.ram01.INIT_04 = 256'h1200B0120113000131B0B012000111011300E001B01300B012000111011300E0,
progmem.ram01.INIT_05 = 256'h00001101130001120101110003110113000112010117000013FF001201130001,
progmem.ram01.INIT_06 = 256'h0001120001110112010111011701130001120001110101110113000112010111,
progmem.ram01.INIT_07 = 256'h02110101110101110113002E01004100001A01011101011101011100001A0113,
progmem.ram01.INIT_08 = 256'h00001A010211001B000011021300011201021101021101021101021101021101,
progmem.ram01.INIT_09 = 256'h01021100001A02021100001202021100001201021100001A0213000212010211,
progmem.ram01.INIT_0A = 256'hFF11010211010211021701021102001202130002120102110000110213000212,
progmem.ram01.INIT_0B = 256'h1102130002120202110102110020110213002E020000112E0200001102001300,
progmem.ram01.INIT_0C = 256'h004100001A031300E0030016030311031300E003001203130002120203110203,
progmem.ram01.INIT_0D = 256'h0303110303110303110000110313000312010311010311000016000317010311,
progmem.ram01.INIT_0E = 256'h030311030311000011031300031200001A030311030311030311030311030311,
progmem.ram01.INIT_0F = 256'h114B0000001A0303110313000312030311030311030311030311030311030311,
progmem.ram01.INIT_10 = 256'h001A0304110413000412000012030411000012030411041300031200001A0304,
progmem.ram01.INIT_11 = 256'h041300E00400130000001104130004120404110413000412040411E004041700,
progmem.ram01.INIT_12 = 256'h0004120204110104110304110417030411020411000011040411000011000411,
progmem.ram01.INIT_13 = 256'h1300041202041101041103041104170304110204110404110000110004110413,
progmem.ram01.INIT_14 = 256'h0004120205110105110405110517030511020511001304051100001100051104,
progmem.ram01.INIT_15 = 256'h1202051101051103051105170305110205113000000013020000110005110513,
progmem.ram01.INIT_16 = 256'h0512020511010511030511051703051102051104051100001100051105130005,
progmem.ram01.INIT_17 = 256'h0000130505110000110005110505110513000500112E05400517000511051300,
progmem.ram01.INIT_18 = 256'h0611000011000611061300051202061101061103061106170306110206113000,
progmem.ram01.INIT_19 = 256'h11061300061200001A0613000612020611010611040611061703061102061104,
progmem.ram01.INIT_1A = 256'h00E006001A061300E0060016060611061300061200001A061300E00600160606,
progmem.ram01.INIT_1B = 256'h1101061101061101061101061101061101061101061106130006124000120613,
progmem.ram01.INIT_1C = 256'h1106071106071106071106071106071106071107130006120107110107110107,
progmem.ram01.INIT_1D = 256'h2E07000011071300071207071101071101071100071107130007120607110607,
progmem.ram01.INIT_1E = 256'h07071107170607112E0700801107071107170307110507110712070012071300,
progmem.ram01.INIT_1F = 256'h0811000011071300E0070013000000110713002E07000211071300071200A011,
progmem.ram01.INIT_20 = 256'hE01107081108170608112E080080110708110817030811060811081300071207,
progmem.ram01.INIT_21 = 256'h11081700081108120800120813000812070811081207081108170608112E0800,
progmem.ram01.INIT_22 = 256'h0811081300081204081108120508110817000012081300081208081108120708,
progmem.ram01.INIT_23 = 256'h0911080811010811081208001208130008122E08008011070811081703081108,
progmem.ram01.INIT_24 = 256'h000009170009112E0800981107091109170009112E0800981109001500091706,
progmem.ram01.INIT_25 = 256'h0609110912090012091300081200981107091109170609110809170609110831,
progmem.ram01.INIT_26 = 256'h0609110913000912000C1107091109170609112E090080110709110917030911,
progmem.ram01.INIT_27 = 256'h2E090080110709110A1703091104091109120900120913000900112E09000917,
progmem.ram01.INIT_28 = 256'h110A17060A112E0A008011070A110A17030A11040A110A1300E0090013090A11,
progmem.ram01.INIT_29 = 256'h0A11090A110A0A110A17010A11070A110013000000110A13000A1200FF11070A,
progmem.ram01.INIT_2A = 256'h0000120000110A00120A13002E0A000011070A110A12070A11080A11080A1109,
progmem.ram01.INIT_2B = 256'h0A001300001200001400230000120A13000A120A0A1100130A13000A120A0013,
progmem.ram01.INIT_2C = 256'h0B110B0B110B0B110B0B110B13000B120A0B110A0B110A0B110A0B110B1300E0,
progmem.ram01.INIT_2D = 256'hB013FFB0120B1300E00B001600B0120B13000B120B0B1100D3110B13000B120B,
progmem.ram01.INIT_2E = 256'h13000B120B1E000B110B170B0B110B1300E00BB01300B0120B0B110B1300E00B,
progmem.ram01.INIT_2F = 256'h110B13000B123C1E0A0B110B0B110B13000B120B0B110B0B110000110B0B110B,
progmem.ram01.INIT_30 = 256'h170B0C110C13000B120B0C110B0C11000C1100AA110C0416000C170B0C11000C,
progmem.ram01.INIT_31 = 256'h0C110B0C110000110B0C110C13000C120B0C110C1EC0FF1600C01B00C013000C,
progmem.ram01.INIT_32 = 256'h0B0C11000C113000CC0C17000C170B0C110A0C110A0C110B0C110C13000C120C,
progmem.ram01.INIT_33 = 256'h00000000000000000C120B0C11000C110C170B0C110A0C110C13000C120B0C11,
progmem.ram01.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
