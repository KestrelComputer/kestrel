`timescale 1ns / 1ps
module NEXYS2(
	output	[2:0]	N2_RED_O,
	output	[2:0]	N2_GRN_O,
	output	[2:1]	N2_BLU_O,
	output			N2_HSYNC_O,
	output			N2_VSYNC_O,
	output			N2_AN0n_O,
	output			N2_AN1n_O,
	output			N2_AN2n_O,
	output			N2_AN3n_O,
	output			N2_CAn_O,
	output			N2_CBn_O,
	output			N2_CCn_O,
	output			N2_CDn_O,
	output			N2_CEn_O,
	output			N2_CFn_O,
	output			N2_CGn_O,
	output			N2_CDPn_O,

	input				N2_50MHZ_I,
	input				N2_BTN0_I,
	input				N2_PS2CLK_I,
	input				N2_PS2DAT_IO,
	
	// SD Card Interface
	output			N2_SD_CLK_O,
	output			N2_SD_MOSI_O,
	output			N2_SD_CS_O,
	output			N2_SD_LED_O,

	input				N2_SD_MISO_I,
	input				N2_SD_WP_I,
	input				N2_SD_CD_I
);

	reg an0n, an1n, an2n, an3n, can, cbn, ccn, cdn, cen, cfn, cgn, cdpn;
	assign N2_AN0n_O = an0n;
	assign N2_AN1n_O = an1n;
	assign N2_AN2n_O = an2n;
	assign N2_AN3n_O = an3n;
	assign N2_CAn_O  = can;
	assign N2_CBn_O  = cbn;
	assign N2_CCn_O  = ccn;
	assign N2_CDn_O  = cdn;
	assign N2_CEn_O  = cen;
	assign N2_CFn_O  = cfn;
	assign N2_CGn_O  = cgn;
	assign N2_CDPn_O = cdpn;

	wire	[15:1]	cpu_adr_o;
	wire				cpu_we_o;
	wire				cpu_cyc_o;
	wire				cpu_stb_o;
	wire	[1:0]		cpu_sel_o;
	wire	[15:0]	cpu_dat_o;
	wire				cpu_ack_i;
	wire	[15:0]	cpu_dat_i;

	wire				kia_ack_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_stb_i;

	wire				gpia_ack_o;
	wire	[15:0]	gpia_dat_o;
	wire				gpia_stb_i;
	wire	[15:0]	gpia_port_o;

	assign N2_SD_CLK_O	= gpia_port_o[3];
	assign N2_SD_MOSI_O	= gpia_port_o[2];
	assign N2_SD_CS_O		= gpia_port_o[1];
	assign N2_SD_LED_O	= gpia_port_o[0];

	wire				progmem_ack_o;
	wire	[15:0]	progmem_dat_o;
	wire				progmem_stb_i;

	wire				vidmem_ack_o;
	wire	[15:0]	vidmem_dat_o;
	wire				vidmem_stb_i;

	wire				mgia_25mhz_o;
	wire	[13:1]	mgia_adr_o;
	wire				mgia_cyc_o;
	wire				mgia_stb_o;
	wire	[15:0]	mgia_dat_i;
	wire				mgia_ack_i;

	wire				cpu_bus_cycle;
	wire				no_peripheral_addressed;

	assign cpu_bus_cycle 				= cpu_cyc_o & cpu_stb_o;
	assign progmem_stb_i 				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b00);		// 0000-3FFF : Program Memory
	assign kia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB00);		// B000-B003 : KIA
	assign gpia_stb_i						= cpu_bus_cycle & (cpu_adr_o[15:4] == 12'hB01);		// B010-B013 : GPIA 
	assign vidmem_stb_i  				= cpu_bus_cycle & (cpu_adr_o[15:14] == 2'b11);		// C000-FFFF : Video Memory
	assign no_peripheral_addressed 	= (~progmem_stb_i & ~kia_stb_i & ~vidmem_stb_i & ~gpia_stb_i);

	wire	[15:0]	progmem_mask 		= {16{progmem_stb_i}};
	wire	[7:0]		kia_mask				= {8{kia_stb_i}};
	wire	[15:0]	vidmem_mask			= {16{vidmem_stb_i}};
	wire	[15:0]	gpia_mask			= {16{gpia_stb_i}};
	assign			cpu_dat_i			= (progmem_mask & progmem_dat_o) | (vidmem_mask & vidmem_dat_o) | {8'b00000000, (kia_mask & kia_dat_o)} | (gpia_mask & gpia_dat_o);
	assign			cpu_ack_i			= (progmem_stb_i & progmem_ack_o) | (vidmem_stb_i & vidmem_ack_o) | (kia_stb_i & kia_ack_o) | (gpia_stb_i & gpia_ack_o) | no_peripheral_addressed;

	always begin
		an0n <= 1'b1;
		an1n <= 1'b1;
		an2n <= 1'b1;
		an3n <= 1'b1;
		can  <= 1'b1;
		cbn  <= 1'b1;
		ccn  <= 1'b1;
		cdn  <= 1'b1;
		cen  <= 1'b1;
		cfn  <= 1'b1;
		cgn  <= 1'b1;
		cdpn <= 1'b1;
	end
	
	S16X4 cpu(
		.adr_o(cpu_adr_o),
		.we_o (cpu_we_o),
		.cyc_o(cpu_cyc_o),
		.stb_o(cpu_stb_o),
		.sel_o(cpu_sel_o),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i),
		.clk_i(mgia_25mhz_o),
		.res_i(N2_BTN0_I)
	);
	
	KIA kia(
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o),
		.CLK_I(mgia_25mhz_o),
		.RES_I(N2_BTN0_I),
		.ADR_I(cpu_adr_o[1]),
		.WE_I (cpu_we_o),
		.CYC_I(cpu_cyc_o),
		.STB_I(kia_stb_i),

		.D_I  (N2_PS2DAT_IO),
		.C_I  (N2_PS2CLK_I)
	);

	GPIA gpia(
		.RST_I(N2_BTN0_I),
		.CLK_I(mgia_25mhz_o),
		.ADR_I(cpu_adr_o[1]),
		.CYC_I(cpu_cyc_o),
		.STB_I(gpia_stb_i),
		.WE_I(cpu_we_o),
		.DAT_I(cpu_dat_o),
		.DAT_O(gpia_dat_o),
		.ACK_O(gpia_ack_o),
		.PORT_I({13'h0000, N2_SD_MISO_I, N2_SD_WP_I, N2_SD_CD_I}),
		.PORT_O(gpia_port_o)
	);

	VRAM16K progmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(progmem_ack_o),
		.A_DAT_O(progmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(progmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ADR_I(13'b1111111111111),
		.B_CYC_I(1'b1),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(1'b0),
		.B_WE_I (1'b1)
	);

	VRAM16K vidmem(
		.CLK_I  (mgia_25mhz_o),

		.A_ACK_O(vidmem_ack_o),
		.A_DAT_O(vidmem_dat_o),
		.A_ADR_I(cpu_adr_o[13:1]),
		.A_CYC_I(cpu_cyc_o),
		.A_DAT_I(cpu_dat_o),
		.A_SEL_I(cpu_sel_o),
		.A_STB_I(vidmem_stb_i),
		.A_WE_I (cpu_we_o),

		.B_ACK_O(mgia_ack_i),
		.B_DAT_O(mgia_dat_i),
		.B_ADR_I(mgia_adr_o[13:1]),
		.B_CYC_I(mgia_cyc_o),
		.B_DAT_I(16'hFFFF),
		.B_SEL_I(2'b11),
		.B_STB_I(mgia_stb_o),
		.B_WE_I (1'b0)
	);

	MGIA mgia(
		.HSYNC_O			(N2_HSYNC_O),
		.VSYNC_O			(N2_VSYNC_O),
		.RED_O			(N2_RED_O),
		.GRN_O			(N2_GRN_O),
		.BLU_O			(N2_BLU_O),
		.MGIA_ADR_O		(mgia_adr_o[13:1]),
		.MGIA_CYC_O		(mgia_cyc_o),
		.MGIA_STB_O		(mgia_stb_o),
		.CLK_O_25MHZ	(mgia_25mhz_o),
		.CLK_I_50MHZ	(N2_50MHZ_I),
		.RST_I			(N2_BTN0_I),
		.MGIA_DAT_I		(mgia_dat_i),
		.MGIA_ACK_I		(mgia_ack_i)
	);
	
defparam
progmem.ram00.INIT_00 = 256'h03FFFF0B0B0B0B0BF303030303ABABAB03FF0000000000000000220044008200,
progmem.ram00.INIT_01 = 256'h00006CE00310156C00005CE00D10155C0000FF6BCB8BCB6BF303030303ABABAB,
progmem.ram00.INIT_02 = 256'h00B4E0B40000AAE0AA0000A0E0A0000096E09600008CE08C0000007C16FF317C,
progmem.ram00.INIT_03 = 256'h00F2002EF2000000DE0112D4EAE0DE0000D2012ED20000C8E0C80000BEE0BE00,
progmem.ram00.INIT_04 = 256'h12F7121532000022E004101522000016002E1600000A002E0A0000FE012EFE00,
progmem.ram00.INIT_05 = 256'h6E12120812166E0000005A1212FD12155A000000461212FB1215460000003212,
progmem.ram00.INIT_06 = 256'h12FF1414B200009C2E1212615CA8E09C000000821212041216488EE082000000,
progmem.ram00.INIT_07 = 256'hFA0000E4E0D0F6E070F0E0E40000CEE0B4E0E0146430CE0000B2E0B8CA1E1414,
progmem.ram00.INIT_08 = 256'hFAE0E63CE0E636E0E630E0E62AE0E624E0E61EE0E618E0E612E0E60CE0E606E0,
progmem.ram00.INIT_09 = 256'h7A000040E0FC76E0FC70E0FC6AE0FC64E0FC5EE0FC58E0FC52E0FC4CE0400000,
progmem.ram00.INIT_0A = 256'hC2E0ACE0BC0E17AC0000009C0E01319C00007AE04298E09E92E0848CE03486E0,
progmem.ram00.INIT_0B = 256'hFA000000EA120031EA0000ACE09EE6E0E60000DCE0ACE09ED2E0D6000CC8E0B6,
progmem.ram00.INIT_0C = 256'h42E046000C38E0CA32E026000010E0EC22E010043010000000FA121201100831,
progmem.ram00.INIT_0D = 256'h1778000026E01274E026E0FC6AE06E001860E026E09E56E05A00004CE026E09E,
progmem.ram00.INIT_0E = 256'hA6E0C0BCE0C000011016A6000078E028A2E078E0EC98E09C006E8EE078E0880E,
progmem.ram00.INIT_0F = 256'hE0EEE0FE0E17EE0000CAE0CAE09EE6E0EA000CDCE0A8D6E0CA0000A6E0A2C6E0,
progmem.ram00.INIT_10 = 256'hE040E0F4E010013A116E2EE0EEE09E24E028005E1AE03A00F410E0CC0AE08E04,
progmem.ram00.INIT_11 = 256'h9E80E084000C76E0CA70E05AE06A0E175A0000EEE09E56E05600004CE0F4461E,
progmem.ram00.INIT_12 = 256'hC40E17B40000980C2E009803AE11F4A4E09800005AE09E94E09400F48AE05AE0,
progmem.ram00.INIT_13 = 256'h000CFEE098F8E0EC000000B410129AE4E0B4E09EDAE0DE000CD0E0ACCAE0B4E0,
progmem.ram00.INIT_14 = 256'h00243EE07C38E00E0000100031200000ECE09E1CE01C00D412E0ECE09E08E00C,
progmem.ram00.INIT_15 = 256'h7A000000200EFF319E70E020E0AE66E07A60E0F05AE05C54E0B64EE0EE48E06A,
progmem.ram00.INIT_16 = 256'h18121A1821B000009CE07CACE01A009C00007AE0801A1E021A141A0023981A17,
progmem.ram00.INIT_17 = 256'h02E0F60000D4E0B2F2E0B2ECE0B2E6E0B2E0E0D4000000B01A12501A14180213,
progmem.ram00.INIT_18 = 256'h2E01120110152E000018E0F82AE01A3630180000F6E0D614E0D60EE0D608E0D6,
progmem.ram00.INIT_19 = 256'h8600307CE070000000561212FE12164462E05600000042121201121542000000,
progmem.ram00.INIT_1A = 256'hC2E044BCE0B000008EE072ACE01AA6E0181C30449AE08E000070E076000486E0,
progmem.ram00.INIT_1B = 256'h00CAE090FAE0B2F4E008EEE0EE001716F41230DCE07ED6E0CA0000B0E000009E,
progmem.ram00.INIT_1C = 256'hE0003EE01A38E0183C30442CE0200000FEE0901CE004001E0E1612300AE0FE00,
progmem.ram00.INIT_1D = 256'h42E0907CE0CC76E00870E070000E76123060E0225AE09E54E0584EE042000020,
progmem.ram00.INIT_1E = 256'h85FFFFB51FFFFFF1FF62FFF10080E090A2E0049CE09C003092E09E8CE0800000,
progmem.ram00.INIT_1F = 256'hDF77BB97FDC5EF7BF5B7FDDF7FAF7BEFEDEBFBF7F7DDEDF85FBFFFFFFF5FFC2F,
progmem.ram00.INIT_20 = 256'h9249247C97F9BFCBEC7B2FF8BFE2FBFFFF7717EE7FFFFFF8F71749775FB9F75F,
progmem.ram00.INIT_21 = 256'h0000000000000000000000000000000000000000005E2FFFAECA57DFFD544524,
progmem.ram00.INIT_22 = 256'hF7E5BFDFBBDBCB7BDDBBBFBFFB44F8FFF9FF2FF2F92400000000000000000000,
progmem.ram00.INIT_23 = 256'hFEB777EE2DFFFFFFFFFFFF5FFF2F7DDDDFEFF7FFFFE5FCFFBEBF2FEEEFDBDF65,
progmem.ram00.INIT_24 = 256'hFFEFFFFFE2FEFEFFFBF8FFF5BFFFFFFF8BFEFFFF498BFFE26F8924792E7BEDFB,
progmem.ram00.INIT_25 = 256'hBFE5CBFFFF97EFFF2FFFFFFFBF77EFF7EEFFC9E2577DFFDEFFC5F1FFFF7FFFF7,
progmem.ram00.INIT_26 = 256'hF7FCFFEFEFEFBEFB8BF7FFFFEFF897FFFFFFFFEFFFF6DFFFF6FBCAF7FF7FFF57,
progmem.ram00.INIT_27 = 256'h5FBCCAAF2FCBDFF8BF2CBEBF2F0BFFDFFFF6FFEFBAC5FF00000400107FEEFFFF,
progmem.ram00.INIT_28 = 256'hFFFE5B7F2FDF7E5F17EFFE78F9EFBB2BB9F7FFFFFFC5FFFF491222912489F9EE,
progmem.ram00.INIT_29 = 256'hFCDD17DFBF0A16E0807F24EF2BFCFCFFFFFEF2FDEFF67FBFBE77FDEE775EBFDD,
progmem.ram00.INIT_2A = 256'h492492492492492448F217C5FE77DFFFFE3BF7DFBFFFFDC5F77FDFBFDF775DFB,
progmem.ram00.INIT_2B = 256'h4992644924669992269249FFF75FFFFF22E8FDAFF2FF2F242492492466666692,
progmem.ram00.INIT_2C = 256'h4999922664249264996699264992494999922664242664494924266449492426,
progmem.ram00.INIT_2D = 256'hFF1FEFFFE5AFFEDFD7EF88F8AF32DC7FDF644999922664249292266449999249,
progmem.ram00.INIT_2E = 256'hDF7FADFDDFFFFF17FFFFCAFFFFF9FFFFDEFFFFFC24AFFFE5FF494491FE2EDFFF,
progmem.ram00.INIT_2F = 256'hCBF2F1D9FEFB5F78FF7FFBFFC6F67FFFFF090000000000000020894989922497,
progmem.ram00.INIT_30 = 256'h0000000000000000EFFFF1EFF7BEDFF7FDF7BECB3BFD7777777DFFE5EE972292,
progmem.ram00.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram00.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

defparam
progmem.ram01.INIT_00 = 256'h180FFFD0D0D0D0D0CFC0C0C8C8CA6232180F0000000000000000071E071E071E,
progmem.ram01.INIT_01 = 256'h130000120000120013000012000012001300FFD6D3D1D3D6CFC0C0C8C8CA6232,
progmem.ram01.INIT_02 = 256'h00001200130000120013000012001300001200130000120013002E0000031100,
progmem.ram01.INIT_03 = 256'h00000011001300E0000016000011001300000011001300001200130000120013,
progmem.ram01.INIT_04 = 256'h13FFB012011300011200B0120113000100110113000100110113000000110013,
progmem.ram01.INIT_05 = 256'h01B01300B012011300E001B013FFB012011300E001B013FFB012011300E001B0,
progmem.ram01.INIT_06 = 256'h13FF00120113000131B0B012010111011300E001B01300B012010111011300E0,
progmem.ram01.INIT_07 = 256'h0113000112010111010111011300011201011100001101130001120101170000,
progmem.ram01.INIT_08 = 256'h0112010211010211010211010211010211010211010211010211010211010211,
progmem.ram01.INIT_09 = 256'h0213000212010211010211010211010211010211010211010211010211021300,
progmem.ram01.INIT_0A = 256'h021102120200120213002E020000110213000212020211010211010211010211,
progmem.ram01.INIT_0B = 256'h0213002E02000211021300021202021102170102110212020211021701021100,
progmem.ram01.INIT_0C = 256'h031103170103110003110313000312020311000011031300E002001300000011,
progmem.ram01.INIT_0D = 256'h1203130003120303110312020311031701031103120203110317010311031202,
progmem.ram01.INIT_0E = 256'h0312000311031700001203130003120303110312020311031700031103120300,
progmem.ram01.INIT_0F = 256'h1103120300120313000312031202031103170103110303110313000312000311,
progmem.ram01.INIT_10 = 256'h0004110331000004170004110312020411041700041104170004110304110004,
progmem.ram01.INIT_11 = 256'h0204110417010411000411041204001204130003120204110417010411030417,
progmem.ram01.INIT_12 = 256'h0400120413000400112E04000417000411041300041202041104170004110412,
progmem.ram01.INIT_13 = 256'h17010411000411041300E0040013040411041202041104170104110004110412,
progmem.ram01.INIT_14 = 256'h1701051102051100130000001105130004120205110517000511041202051105,
progmem.ram01.INIT_15 = 256'h0513002E05000011020511051202051103051103051104051104051104051105,
progmem.ram01.INIT_16 = 256'h0023000012051300051205051100130513000512050013000012000011050012,
progmem.ram01.INIT_17 = 256'h06110513000512050511050511050511050511051300E0050013000012000014,
progmem.ram01.INIT_18 = 256'h06001600B012061300061205061100D311061300051205061105061105061105,
progmem.ram01.INIT_19 = 256'h0617060611061300E006B013FFB012060611061300E006B01300B012061300E0,
progmem.ram01.INIT_1A = 256'h061106061106130006120606110606110000110606110613000612061E000611,
progmem.ram01.INIT_1B = 256'h00061206061106061100061106041600061706061100061106130006123C1E05,
progmem.ram01.INIT_1C = 256'h12070711060711000011060711071300061206071107C0130007170607110613,
progmem.ram01.INIT_1D = 256'h0712060711060711000711071700071706071105071105071106071107130007,
progmem.ram01.INIT_1E = 256'hFE17FFBFF8FE9F5FFFF7FF7F0007120607110007110717060711050711071300,
progmem.ram01.INIT_1F = 256'hFDDFEFE5FFFBBF16F5FF5EBFFFD5D55DBAEFDFDEEBAFEFBFFFBCFCFFFFFFBC0B,
progmem.ram01.INIT_20 = 256'h492492BFF97FCBFCBFFF99BFFFFC17FF8BFFF1FFEEC5BBBF7FFF33F2EF71F8FB,
progmem.ram01.INIT_21 = 256'h0000000000000000000000000000000000000000004077EFF2FCDDF6EF975592,
progmem.ram01.INIT_22 = 256'hF9F2FFFDEFFDFFBFFB7FF7FC5F9722977FFFFF497DBF01000000000000000000,
progmem.ram01.INIT_23 = 256'h2E7FFBFFDFFEFFFFFFFF85FFF9FFBCF7777DDD62FBF25F17FBDBFDFFEDFEBDFF,
progmem.ram01.INIT_24 = 256'hCBF7FF9725FF2FFF2FBFFFFFDFD8FF8BF25FFFE222161DCEBF11887F5BBFF9BC,
progmem.ram01.INIT_25 = 256'hF6FFFFFFFFFFFDFFFFFFE5CB8BB8BF7EFBDF17DF7FFCFF2BFFFF57FFFFFFF1FF,
progmem.ram01.INIT_26 = 256'hFF5FFFFFFBBFFBEFBEFDFFFFFFBEFFFFFF62FF2FE22F65E257BFFF7E2FFFD9FF,
progmem.ram01.INIT_27 = 256'hF8BCF22BFC89BF5F7758EEBBF8FCFBFF0B17FFDDFFDE2F1200400000BFF1EEFF,
progmem.ram01.INIT_28 = 256'h5FDFBFFEC5BF2FBFBCDFB7BB7F778BF37EEFFBFEFF8BEFFF8A24491148127FF1,
progmem.ram01.INIT_29 = 256'h0FF77FEFDFBF0B7EF9C749F7BEBEBFCBCB77EF8BF6B5F7EBFBD7DEFB9649F6FF,
progmem.ram01.INIT_2A = 256'h249249249249249291FCCBFF2FFFBBFFCAFFFFBFFFE08BFFF8FD17C578FFF1F8,
progmem.ram01.INIT_2B = 256'h9966992692492664494924C6FFFFECFF22B1FFFEFCFFFE4C9249249249666666,
progmem.ram01.INIT_2C = 256'h9226644999924999264992649966249226644999924999922692499992269249,
progmem.ram01.INIT_2D = 256'hFFFFFFEFFF7EF7FFD7D725BFFFC55FE22F859226644999924964499992266424,
progmem.ram01.INIT_2E = 256'hDFDDFFFFEB7777CBCBFFF7FFFF7FFF2FFFFFFFBFB292FC7FFF2592225CFDFFEF,
progmem.ram01.INIT_2F = 256'hF7F7FB7FDFFEFEFCDF7FD97D5F2F7EDF176200000000000000001224244448DE,
progmem.ram01.INIT_30 = 256'h00000000000000007EBD6F75FE5FFBFFFFCB5FFBFFEFBBF7FFFFFFE55EE54449,
progmem.ram01.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
progmem.ram01.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
